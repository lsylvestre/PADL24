library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 11);
       signal result : out value(0 to 57));
       
end entity;
architecture rtl of main is

  type t_state is (compute1859);
  signal state: t_state;
  type t_state_var5313 is (compute2976, pause_setI2977, pause_setI2978, pause_setI2979, pause_setI2980, pause_setI2981, pause_setI2982, pause_setI2983, pause_setI2984, pause_setI2985, pause_setI2986, pause_setI2987, pause_setI2988, pause_setI2989, pause_setI2990, pause_setI2991, pause_setI2992, pause_setI2993, pause_setI2994, pause_setI2995, pause_setI2996, pause_setI2997, pause_setI2998, pause_setI2999, pause_setI3000, pause_setI3001, pause_setI3002, pause_setI3003, pause_setI3004, pause_setI3005, pause_setI3006, pause_setI3007, pause_setI3008, pause_setI3009, pause_setI3010, pause_setI3011, pause_setI3012, pause_setI3013, pause_setI3014, pause_setI3015, pause_setI3016, pause_setI3017, pause_setI3018, pause_setI3019, pause_setI3020, pause_setI3021, pause_setI3022, pause_setI3023, pause_setI3024, pause_setI3025, pause_setI3026, pause_setI3027, pause_setI3028, pause_setI3029, pause_setI3030, pause_setI3031, pause_setI3032, pause_setI3033, pause_setI3034, pause_setI3035, pause_setI3036, pause_setI3037, pause_setI3038, pause_setI3039, pause_setI3040, pause_setI3041, pause_setI3042, pause_setI3043, pause_setI3044, pause_setI3045, pause_setI3046, pause_setI3047, pause_setI3048, pause_setI3049, pause_setI3050, pause_setI3051, pause_setI3052, pause_setI3053, pause_setI3054, pause_setI3055, pause_setI3056, pause_setI3057, pause_setI3058, pause_setI3059, pause_setI3060, pause_setI3061, pause_setI3062, pause_setI3063, pause_setI3064, pause_setI3065, pause_setI3066, pause_setI3067, pause_setI3068, pause_setI3069, pause_setI3070, pause_setI3071, pause_setI3072, pause_setI3073, pause_setI3074, pause_setI3075, pause_setI3076, pause_setI3077, pause_setI3078, pause_setI3079, pause_setI3080, pause_setI3081, pause_setI3082, pause_setI3083, pause_setI3084, pause_setI3085, pause_setI3086, pause_setI3087, pause_setI3088, pause_setI3089, pause_setI3090, pause_setI3091, pause_setI3092, pause_setI3093, pause_setI3094, pause_setI3095, pause_setI3096, pause_setI3097, pause_setI3098, pause_setI3099, pause_setI3100, pause_setI3101, pause_setI3102, pause_setI3103, pause_setI3104, pause_setI3105, pause_setI3106, pause_setI3107, pause_setI3108, pause_setI3109, pause_setI3110, pause_setI3111, pause_setI3112, pause_setI3113, pause_setI3114, pause_setI3115, pause_setI3116, pause_setI3117, pause_setI3118, pause_setI3119, pause_setI3120, pause_setI3121, pause_setI3122, pause_setI3123, pause_setI3124, pause_setI3125, pause_setI3126, pause_setI3127, pause_setI3128, pause_setI3129, pause_setI3130, pause_setI3131, pause_setI3132, pause_setI3133, pause_setI3134, pause_setI3135, pause_setI3136, pause_setI3137, pause_setI3138, pause_setI3139, pause_setI3140, pause_setI3141, pause_setI3142, pause_setI3143, pause_setI3144, pause_setI3145, pause_setI3146, pause_setI3147, pause_setI3148, pause_setI3149, pause_setI3150, pause_setI3151, pause_setI3152, pause_setI3153, pause_setI3154, pause_setI3155, pause_setI3156, pause_setI3157, pause_setI3158, pause_setI3159, pause_setI3160, pause_setI3161, pause_setI3162, pause_setI3163, pause_setI3164, pause_setI3165, pause_setI3166, pause_setI3167, pause_setI3168, pause_setI3169, pause_setI3170, pause_setI3171, pause_setI3172, pause_setI3173, pause_setI3174, pause_setI3175, pause_setI3176, pause_setI3177, pause_setI3178, pause_setI3179, pause_setI3180, pause_setI3181, pause_setI3182, pause_setI3183, pause_setI3184, pause_setI3185, pause_setI3186, pause_setI3187, pause_setI3188, pause_setI3189, pause_setI3190, pause_setI3191, pause_setI3192, pause_setI3193, pause_setI3194, pause_setI3195, pause_setI3196, pause_setI3197, pause_setI3198, pause_setI3199, pause_setI3200, pause_setI3201, pause_setI3202, pause_setI3203, pause_setI3204, pause_setI3205, pause_setI3206, pause_setI3207, pause_setI3208, pause_setI3209, pause_setI3210, pause_setI3211, pause_setI3212, pause_setI3213, pause_setI3214, pause_setI3215, pause_setI3216, pause_setI3217, pause_setI3218, pause_setI3219, pause_setI3220, pause_setI3221, pause_setI3222, pause_setI3223, pause_setI3224, pause_setI3225, pause_setI3226, pause_setI3227, pause_setI3228, pause_setI3229, pause_setI3230, pause_setI3231, pause_setI3232, pause_setI3233, pause_setI3234, pause_setI3235, pause_setI3236, pause_setI3237, pause_setI3238, pause_setI3239, pause_setI3240, pause_setI3241, pause_setI3242, pause_setI3243, pause_setI3244, pause_setI3245, pause_setI3246, pause_setI3247, pause_setI3248, pause_setI3249, pause_setI3250, pause_setI3251, pause_setI3252, pause_setI3253, pause_setI3254, pause_setI3255, pause_setI3256, pause_setI3257, pause_setI3258, pause_setI3259, pause_setI3260, pause_setI3261, pause_setI3262, pause_setI3263, pause_setI3264, pause_setI3265, pause_setI3266, pause_setI3267, pause_setI3268, pause_setI3269, pause_setI3270, pause_setI3271, pause_setI3272, pause_setI3273, pause_setI3274, pause_setI3275, pause_setI3276, pause_setI3277, pause_setI3278, pause_setI3279, pause_setI3280, pause_setI3281, pause_setI3282, pause_setI3283, pause_setI3284, pause_setI3285, pause_setI3286, pause_setI3287, pause_setI3288, pause_setI3289, pause_setI3290, pause_setI3291, pause_setI3292, pause_setI3293, pause_setI3294, pause_setI3295, pause_setI3296, pause_setI3297, pause_setI3298, pause_setI3299, pause_setI3300, pause_setI3301, pause_setI3302, pause_setI3303, pause_setI3304, pause_setI3305, pause_setI3306, pause_setI3307, pause_setI3308, pause_setI3309, pause_setI3310, pause_setI3311, pause_setI3312, pause_setI3313, pause_setI3314, pause_setI3315, pause_setI3316, pause_setI3317, pause_setI3318, pause_setI3319, pause_setI3320, pause_setI3321, pause_setI3322, pause_setI3323, pause_setI3324, pause_setI3325, pause_setI3326, pause_setI3327, pause_setI3328, pause_setI3329, pause_setI3330, pause_setI3331, pause_setI3332, pause_setI3333, pause_setI3334, pause_setI3335, pause_setI3336, pause_setI3337, pause_setI3338, pause_setI3339, pause_setI3340, pause_setI3341, pause_setI3342, pause_setI3343, pause_setI3344, pause_setI3345, pause_setI3346, pause_setI3347, pause_setI3348, pause_setI3349, pause_setI3350, pause_setI3351, pause_setI3352, pause_setI3353, pause_setI3354, pause_setI3355, pause_setI3356, pause_setI3357, pause_setI3358, pause_setI3359, pause_setI3360, pause_setI3361, pause_setI3362, pause_setI3363, pause_setI3364, pause_setI3365, pause_setI3366, pause_setI3367, pause_setI3368, pause_setI3369, pause_setI3370, pause_setI3371, pause_setI3372, pause_setI3373, pause_setI3374, pause_setI3375, pause_setI3376, pause_setI3377, pause_setI3378, pause_setI3379, pause_setI3380, pause_setI3381, pause_setI3382, pause_setI3383, pause_setI3384, pause_setI3385, pause_setI3386, pause_setI3387, pause_setI3388, pause_setI3389, pause_setI3390, pause_setI3391, pause_setI3392, pause_setI3393, pause_setI3394, pause_setI3395, pause_setI3396, pause_setI3397, pause_setI3398, pause_setI3399, pause_setI3400, pause_setI3401, pause_setI3402, pause_setI3403, pause_setI3404, pause_setI3405, pause_setI3406, pause_setI3407, pause_setI3408, pause_setI3409, pause_setI3410, pause_setI3411, pause_setI3412, pause_setI3413);
  signal state_var5313: t_state_var5313;
  type t_state_var5312 is (compute4920, \$706_loop\, \$707_copy_root_in_ram\, \$708_loop\, \$709_aux\, \$710\, \$711_apply\, \$712_offsetclosure_n\, \$713_binop_int\, \$714_compare\, \$715_binop_compare\, \$716_make_block_n\, \$717_branch_if\, \$718_loop_push\, \$719_compbranch\, \$720_w\, \$721_w\, \$722_fill\, \$723_fill\, \$724_w0\, \$725_w1\, \$726_w3\, pause_getI5049, pause_getI5051, pause_getI5053, pause_getI5055, pause_getI5057, pause_getI5059, pause_getI5061, pause_getI5063, pause_getI5067, pause_getI5070, pause_getI5073, pause_getI5076, pause_getI5079, pause_getI5082, pause_getI5085, pause_getI5088, pause_getI5090, pause_getI5092, pause_getI5094, pause_getI5096, pause_getI5099, pause_getI5102, pause_getI5105, pause_getI5108, pause_getI5110, pause_getI5116, pause_getI5118, pause_getI5120, pause_getI5122, pause_getI5125, pause_getI5128, pause_getI5131, pause_getI5134, pause_getI5136, pause_getI5138, pause_getI5140, pause_getI5143, pause_getI5145, pause_getI5147, pause_getI5149, pause_getI5152, pause_getI5154, pause_getI5156, pause_getI5158, pause_getI5160, pause_getI5162, pause_getI5164, pause_getI5170, pause_getI5172, pause_getI5176, pause_getI5178, pause_getI5184, pause_getI5186, pause_getI5188, pause_getI5190, pause_getI5192, pause_getI5195, pause_getI5197, pause_getI5199, pause_getI5205, pause_getI5207, pause_getI5212, pause_getI5215, pause_getI5217, pause_getI5219, pause_getI5226, pause_getI5230, pause_getI5234, pause_getI5236, pause_getI5240, pause_getI5242, pause_getI5244, pause_getI5248, pause_getI5250, pause_getI5252, pause_getI5254, pause_getI5258, pause_getI5260, pause_getI5262, pause_getI5264, pause_getI5268, pause_getI5270, pause_getI5275, pause_getI5277, pause_getI5279, pause_getI5281, pause_getI5289, pause_getI5292, pause_getI5295, pause_getI5298, pause_getI5301, pause_getII5050, pause_getII5052, pause_getII5054, pause_getII5056, pause_getII5058, pause_getII5060, pause_getII5062, pause_getII5064, pause_getII5068, pause_getII5071, pause_getII5074, pause_getII5077, pause_getII5080, pause_getII5083, pause_getII5086, pause_getII5089, pause_getII5091, pause_getII5093, pause_getII5095, pause_getII5097, pause_getII5100, pause_getII5103, pause_getII5106, pause_getII5109, pause_getII5111, pause_getII5117, pause_getII5119, pause_getII5121, pause_getII5123, pause_getII5126, pause_getII5129, pause_getII5132, pause_getII5135, pause_getII5137, pause_getII5139, pause_getII5141, pause_getII5144, pause_getII5146, pause_getII5148, pause_getII5150, pause_getII5153, pause_getII5155, pause_getII5157, pause_getII5159, pause_getII5161, pause_getII5163, pause_getII5165, pause_getII5171, pause_getII5173, pause_getII5177, pause_getII5179, pause_getII5185, pause_getII5187, pause_getII5189, pause_getII5191, pause_getII5193, pause_getII5196, pause_getII5198, pause_getII5200, pause_getII5206, pause_getII5208, pause_getII5213, pause_getII5216, pause_getII5218, pause_getII5220, pause_getII5227, pause_getII5231, pause_getII5235, pause_getII5237, pause_getII5241, pause_getII5243, pause_getII5245, pause_getII5249, pause_getII5251, pause_getII5253, pause_getII5255, pause_getII5259, pause_getII5261, pause_getII5263, pause_getII5265, pause_getII5269, pause_getII5271, pause_getII5276, pause_getII5278, pause_getII5280, pause_getII5282, pause_getII5290, pause_getII5293, pause_getII5296, pause_getII5299, pause_getII5302, pause_setI5065, pause_setI5066, pause_setI5069, pause_setI5072, pause_setI5075, pause_setI5078, pause_setI5081, pause_setI5084, pause_setI5087, pause_setI5098, pause_setI5101, pause_setI5104, pause_setI5107, pause_setI5112, pause_setI5113, pause_setI5114, pause_setI5115, pause_setI5124, pause_setI5127, pause_setI5130, pause_setI5133, pause_setI5142, pause_setI5151, pause_setI5166, pause_setI5167, pause_setI5168, pause_setI5169, pause_setI5174, pause_setI5175, pause_setI5180, pause_setI5181, pause_setI5182, pause_setI5183, pause_setI5201, pause_setI5202, pause_setI5204, pause_setI5209, pause_setI5210, pause_setI5211, pause_setI5214, pause_setI5222, pause_setI5223, pause_setI5224, pause_setI5225, pause_setI5229, pause_setI5233, pause_setI5239, pause_setI5247, pause_setI5257, pause_setI5266, pause_setI5267, pause_setI5272, pause_setI5273, pause_setI5283, pause_setI5284, pause_setI5285, pause_setI5286, pause_setI5287, pause_getI4922, pause_getII4923, pause_setI4921, pause_getI4929, pause_getI4932, pause_getI4935, pause_getII4930, pause_getII4933, pause_getII4936, pause_setI4925, pause_setI4926, pause_setI4927, pause_setI4928, pause_getI4942, pause_getI4945, pause_getI4948, pause_getII4943, pause_getII4946, pause_getII4949, pause_setI4938, pause_setI4939, pause_setI4940, pause_setI4941, pause_getI4951, pause_getII4952, pause_getI4955, pause_getI4960, pause_getI4963, pause_getI4969, pause_getI4972, pause_getII4956, pause_getII4961, pause_getII4964, pause_getII4970, pause_getII4973, pause_setI4954, pause_setI4957, pause_setI4958, pause_setI4959, pause_setI4966, pause_setI4967, pause_setI4968, pause_getI4977, pause_getI4989, pause_getI4992, pause_getI4995, pause_getII4978, pause_getII4990, pause_getII4993, pause_getII4996, pause_setI4979, pause_setI4981, pause_setI4983, pause_setI4985, pause_setI4986, pause_setI4987, pause_getI5000, pause_getII5001, pause_getI5003, pause_getII5004, pause_getI5006, pause_getI5010, pause_getII5007, pause_getII5011, pause_setI5005, pause_setI5009, pause_setI5013, pause_getI5015, pause_getII5016, pause_getI5019, pause_getII5020, pause_setI5018, pause_getI5023, pause_getII5024, pause_setI5022, pause_getI5027, pause_getII5028, pause_setI5026, pause_getI5031, pause_getII5032, pause_setI5030, pause_getI5035, pause_getII5036, pause_setI5034, pause_getI5039, pause_getII5040, pause_setI5038, pause_getI5043, pause_getII5044, pause_setI5042, pause_setI5045, pause_setI5047);
  signal state_var5312: t_state_var5312;
  type array_value_16 is array (natural range <>) of value(0 to 15);
  type array_value_31 is array (natural range <>) of value(0 to 30);
  type array_value_32 is array (natural range <>) of value(0 to 31);
  signal ram : array_value_32(0 to 16383);
  signal \$ram_value\ : value(0 to 31);
  signal \$ram_ptr\ : natural range 0 to 16383;
  signal \$ram_ptr_write\ : natural range 0 to 16383;
  signal \$ram_write\ : value(0 to 31);
  signal \$ram_write_request\ : std_logic := '0';
  signal global_end : array_value_16(0 to 0);
  signal \$global_end_value\ : value(0 to 15);
  signal \$global_end_ptr\ : natural range 0 to 0;
  signal \$global_end_ptr_write\ : natural range 0 to 0;
  signal \$global_end_write\ : value(0 to 15);
  signal \$global_end_write_request\ : std_logic := '0';
  signal code : array_value_31(0 to 421);
  signal \$code_value\ : value(0 to 30);
  signal \$code_ptr\ : natural range 0 to 421;
  signal \$code_ptr_write\ : natural range 0 to 421;
  signal \$code_write\ : value(0 to 30);
  signal \$code_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                 -- if \$ram_write_request\ = '1' then
                    ram(\$ram_ptr_write\) <= \$ram_write\;
                 -- else
                   \$ram_value\ <= ram(\$ram_ptr\);
                 -- end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                 -- if \$global_end_write_request\ = '1' then
                    global_end(\$global_end_ptr_write\) <= \$global_end_write\;
                 -- else
                   \$global_end_value\ <= global_end(\$global_end_ptr\);
                 -- end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                 -- if \$code_write_request\ = '1' then
                    code(\$code_ptr_write\) <= \$code_write\;
                 -- else
                   \$code_value\ <= code(\$code_ptr\);
                 -- end if;
            end if;
        end process;
    
    process(clk)
      variable \$v1557\, \$v1822\
               : value(0 to 1) := (others => '0');
      variable \$713_binop_int_arg\
               : value(0 to 154) := (others => '0');
      variable \$717_branch_if_arg\
               : value(0 to 138) := (others => '0');
      variable \$707_copy_root_in_ram_arg\, \$v3595\, \$v3547\, \$v3596\, 
               \$724_w0_arg\, \$v3589\, \$710_result\, \$v3600\, \$v3611\
               : value(0 to 95) := (others => '0');
      variable \$714_compare_arg\
               : value(0 to 93) := (others => '0');
      variable \$720_w_arg\, \$718_loop_push_arg\, \$706_loop_arg\, 
               \$721_w_arg\
               : value(0 to 63) := (others => '0');
      variable \$v3633\, \$v3628\, \$v3646\, \$v3654\, \$v3639\
               : value(0 to 32) := (others => '0');
      variable \$v3569\, \$v3566\, \$v3609\, \$v3687\, \$v3651\, \$v3693\, 
               \$v3694\, \$v3695\, \$v3610\, \$v3653\, \$v3427\, \$1101\, 
               \$v3698\, \$v3549\, \$v3629\, \$v3563\, \$v3558\, \$v3545\, 
               \$v3634\, \$v3528\, \$v3637\, \$v3614\, \$v3701\, \$v3689\, 
               \$v3699\, \$v3655\, \$v3697\, \$v3616\, \$v3530\, \$v3691\, 
               \$v3638\, \$v3615\, \$v3681\, \$v3644\, \$v3650\, \$v3608\, 
               \$v3647\, \$v3542\, \$v3486\, \$v3645\, \$v3690\, \$v3683\, 
               \$v3622\, \$v3700\, \$v3640\, \$v3643\, \$v3551\, \$v3652\, 
               \$v3529\, \$v3446\, \$v3632\, \$v3685\, \$v3487\
               : value(0 to 47) := (others => '0');
      variable \$v232\, \$v1814\, \$v1545\, \$v1549\, \$v1820\
               : value(0 to 122) := (others => '0');
      variable \$v5291\, \$547_o\, \$v5294\, \$v5297\, \$v5300\
               : value(0 to 7) := (others => '0');
      variable \$5459_sp\, \$975_sp\, \$1579\, \$803_sp\, \$967\, \$951_sp\, 
               \$722_fill_result\, \$5370_sp\, \$1297_sp\, \$1285_sp\, 
               \$859_sp\, \$1567_next\, \$893_sp\, \$792_sp\, \$5448_sp\, 
               \$5392_sp\, \$883_ofs\, \$1179_sp\, \$1288_sp\, \$1278_sp\, 
               \$5461_sp\, \$720_w_result\, \$1568_next\, \$5397_sp\, 
               \$718_loop_push_result\, \$1243_sp\, \$726_w3_result\, 
               \$879_sp\, \$785_sp\, \$976\, \$1038_sp\, \$708_loop_result\, 
               \$1180_sp\, \$814_sp\, \$1312_sp\, \$5402_sp\, 
               \$707_copy_root_in_ram_result\, \$763_sp\, \$709_aux_result\, 
               \$1305_sp\, \$888_idx\, \$778_sp\, \$901_sp\, \$5434_sp\, 
               \$1620\, \$764_sp\, \$5372_sp\, \$912_sp\, \$5427_sp\, 
               \$923_sp\, \$5557_sp\, \$1332_sp\, \$5387_sp\, \$1284_sp\, 
               \$723_fill_result\, \$936_sp\, \$1565_next\, \$5114\, 
               \$902_sp\, \$724_w0_result\, \$1277_sp\, \$970_sp\, \$875_sp\, 
               \$1275_sp\, \$752_sp\, \$5085\, \$1276_sp\, \$5563_sp\, 
               \$894_sp\, \$1581_next\, \$819_sp\, \$5141\, \$5377_sp\, 
               \$903_sp\, \$762_sp\, \$5566_sp\, \$1566\, \$5382_sp\, 
               \$5463_sp\, \$5441_sp\, \$1139_sp\, \$820_sp\, \$5560_sp\
               : value(0 to 15) := (others => '0');
      variable \$708_loop_arg\
               : value(0 to 111) := (others => '0');
      variable \$710_arg\
               : value(0 to 167) := (others => '0');
      variable result1857
               : value(0 to 57) := (others => '0');
      variable \$716_make_block_n_id\, \$706_loop_id\, \$719_compbranch_id\, 
               \$723_fill_id\, \$710_id\, \$722_fill_id\, 
               \$707_copy_root_in_ram_id\, \$712_offsetclosure_n_id\, 
               \$708_loop_id\, \$726_w3_id\, \$725_w1_id\, \$714_compare_id\, 
               \$711_apply_id\, \$720_w_id\, \$718_loop_push_id\, 
               \$713_binop_int_id\, \$724_w0_id\, \$709_aux_id\, 
               \$715_binop_compare_id\, \$717_branch_if_id\, \$721_w_id\
               : value(0 to 11) := (others => '0');
      variable \$746_argument3\, \$885\, \$740\, \$v5256\, \$1152_arg\, 
               \$v5238\, \$v5246\, \$v5228\, \$745_argument2\, \$1218_res\, 
               \$1055\, \$747\, \$744_argument1\, \$v5232\
               : value(0 to 30) := (others => '0');
      variable \$712_offsetclosure_n_arg\
               : value(0 to 137) := (others => '0');
      variable \$v1809\, \$v1527\, \$v495\
               : value(0 to 10) := (others => '0');
      variable \$725_w1_arg\
               : value(0 to 103) := (others => '0');
      variable \$v1808\
               : value(0 to 9) := (others => '0');
      variable \$716_make_block_n_arg\
               : value(0 to 235) := (others => '0');
      variable \$v3477\, \$1530\, \$v3419\
               : value(0 to 127) := (others => '0');
      variable \$v5309\, \$v2501\, \$v2498\, \$v5021\, \$v2769\, \$v2820\, 
               \$v2534\, \$v2928\, \$v2516\, \$v3428\, \$v2652\, \$v4934\, 
               \$v2868\, \$v2580\, \$v2592\, \$v1556\, \$v2791\, \$v4976\, 
               \$v2748\, \$v5014\, \$v2809\, \$v2774\, \$v3532\, \$v2764\, 
               \$v3417\, \$v2812\, \$v2854\, \$v2762\, \$v2768\, \$v2617\, 
               \$v2505\, \$v5274\, \$v3548\, \$v2783\, \$v3567\, \$v2731\, 
               \$v2520\, \$548_rdy\, \$v5203\, \$v1818\, result4918, 
               \$v2875\, \$v2781\, \$v2653\, \$714_compare_result\, \$v2660\, 
               \$v2788\, \$v2730\, \$v2651\, \$v2646\, \$725_w1_result\, 
               \$v2607\, \$v2726\, \$v5310\, \$v2540\, \$v3416\, \$v3575\, 
               \$v2630\, \$v3441\, \$v4971\, \$v2627\, \$v2670\, \$v3599\, 
               \$v14\, \$v2712\, \$v2931\, \$v5303\, \$v3559\, \$v2545\, 
               \$v2866\, \$v2782\, \$v3606\, \$v2873\, \$v2656\, \$v2581\, 
               \$1127_b\, \$v2818\, \$v3674\, \$v2912\, \$v2897\, \$v2844\, 
               \$v2761\, \$v2513\, \$v2500\, \$v2837\, \$v1556_init\, 
               \$v2800\, \$v3636\, \$v2801\, \$v2691\, \$v3660\, \$v2914\, 
               \$v2564\, \$v2923\, \$v2704\, \$v2508\, \$v2725\, \$v2503\, 
               \$v3457\, \$v2879\, \$v2714\, \$v2542\, \$v2900\, \$v2833\, 
               \$v2700\, \$v2524\, \$v2780\, \$v2523\, \$v2901\, \$v2933\, 
               \$v5307\, \$706_loop_result\, \$v2838\, \$v2688\, \$v3550\, 
               \$v3415\, \$v2894\, \$v2546\, \$v2728\, \$v1557_init\, 
               \$v3617\, \$v2910\, \$v2680\, \$v5046\, \$v2796\, \$v3661\, 
               \$v2706\, \$v2649\, \$v2870\, \$v2635\, \$v3626\, \$v2773\, 
               \$v2543\, \$v3642\, \$v2776\, \$v2566\, \$v2760\, \$v2674\, 
               \$v2707\, \$v2589\, \$v4953\, \$v4931\, \$v3592\, \$v2798\, 
               \$v2789\, \$v2497\, \$v2926\, \$v2790\, \$v2699\, \$v2679\, 
               \$v2594\, \$v2636\, \$v2729\, \$v2766\, \$v2701\, \$v2687\, 
               \$v2664\, \$v2806\, \$v2932\, \$v4980\, \$v2579\, \$v3670\, 
               \$v1549_init\, \$v3665\, \$v1823\, \$v3519\, \$v2573\, 
               \$v2920\, \$v2531\, \$v2514\, \$v2834\, \$v2824\, \$v5025\, 
               \$v2696\, \$v2684\, \$v3631\, \$v2905\, \$v2904\, \$v2517\, 
               \$v2723\, \$v2889\, \$v2795\, \$v5308\, \$v3684\, \$v2869\, 
               \$v3676\, \$v2823\, \$v2530\, \$v2930\, \$v2862\, \$v4998\, 
               \$v5048\, \$v2765\, \$v2686\, \$v2563\, \$v2548\, \$v3458\, 
               \$v2860\, \$v2848\, \$v3649\, \$v2740\, \$v2565\, \$v2626\, 
               \$v3504\, \$v3444\, \$v1860\, \$v4982\, \$v2861\, \$v2705\, 
               \$v4988\, \$v2609\, \$v3503\, \$v2721\, \$v2720\, \$v2908\, 
               \$v2578\, \$v2568\, \$v2927\, \$v3443\, \$v2763\, \$v2711\, 
               \$v2683\, \$v3604\, \$v2676\, \$v4962\, \$v2727\, \$v2872\, 
               \$v2692\, \$v5041\, result2974, \$v2515\, \$v2570\, \$v2867\, 
               \$v2586\, rdy2975, \$v3601\, \$v2681\, \$v2536\, \$v2644\, 
               \$v2596\, \$1196_res\, \$v2575\, \$v2598\, \$v2601\, \$v2518\, 
               \$v2697\, \$v2896\, \$v2832\, \$v2554\, \$v2577\, \$v2917\, 
               \$v2831\, \$v2892\, \$v2841\, \$v2622\, \$v5288\, \$v3625\, 
               \$v2767\, \$v3682\, \$v2510\, \$v5311\, \$v2847\, \$v2591\, 
               \$v3666\, \$v2895\, \$v2799\, \$v2849\, \$v2797\, \$v2843\, 
               \$v2807\, \$v5033\, \$v2645\, \$v2924\, \$v2857\, \$v2620\, 
               \$v2826\, \$v2709\, \$v2794\, \$v2759\, \$v3516\, \$v3672\, 
               \$v1563_init\, \$v2830\, \$v2572\, \$v2708\, \$v3663\, 
               \$v3671\, \$v3535\, \$v2642\, \$v2661\, \$v2643\, \$v2815\, 
               \$v2746\, \$v2903\, \$v2856\, \$v3619\, \$v2913\, \$v3573\, 
               \$v2606\, \$v2504\, \$v2785\, \$v2593\, \$v2551\, \$v2784\, 
               \$v2745\, \$v3478\, \$v2600\, \$v2732\, \$v2561\, \$v2506\, 
               \$v2499\, \$v2718\, \$v2628\, \$v1810\, \$v5037\, \$v2906\, 
               \$v2657\, \$v2667\, \$v2871\, \$v2851\, \$v2717\, \$v2659\, 
               \$v5194\, \$v1825\, \$v2615\, \$v2507\, \$v3620\, \$v2828\, 
               \$v3570\, \$v2777\, \$v2595\, \$v2535\, \$v5012\, \$v2840\, 
               \$v2810\, \$v2529\, \$v2668\, \$v2647\, \$v2571\, \$v3572\, 
               \$v2881\, \$v2878\, \$v3612\, \$v2538\, \$v2537\, \$v2770\, 
               \$v2886\, \$v2698\, \$v2532\, \$v3533\, \$v2880\, \$v2677\, 
               \$v2758\, \$v2613\, \$v1545_init\, \$v2654\, \$v2816\, 
               \$v2863\, \$v2850\, \$v3658\, \$v2576\, \$v2929\, \$v3618\, 
               \$v2755\, \$v2559\, \$v2703\, \$v2666\, \$v2528\, \$v2716\, 
               \$v2814\, \$v2663\, \$v2819\, \$v4997\, \$v2682\, \$v3675\, 
               \$v2621\, \$v2888\, \$v2853\, \$v2771\, \$721_w_result\, 
               \$v2637\, \$v2623\, \$v3576\, \$v2802\, \$v2778\, \$v3447\, 
               \$v2555\, \$v3552\, \$v2859\, \$v2685\, \$v3623\, \$v2738\, 
               \$v2911\, \$v2618\, \$v2552\, \$v4984\, \$v2512\, \$v2925\, 
               \$v3668\, \$v2672\, \$v3593\, \$v3460\, \$v2821\, \$v3696\, 
               \$v2736\, \$v2616\, \$v2648\, \$v2629\, \$v3506\, \$v2915\, 
               \$v2724\, \$v3564\, \$v2902\, \$v2662\, \$v2753\, \$v2855\, 
               \$v2665\, \$v2852\, \$v2619\, \$v3704\, \$v2918\, \$v2742\, 
               \$v2839\, \$v2813\, \$v3673\, \$v2749\, \$v3594\, 
               \$v3419_init\, \$v3657\, \$v2793\, \$v2671\, \$v2560\, 
               \$v2527\, \$v3591\, \$v3505\, \$v2590\, \$v4965\, \$v3597\, 
               \$v3692\, \$v5304\, \$v2673\, rdy4919, \$v2715\, \$v2584\, 
               \$v2690\, \$v2611\, \$v2864\, \$v3669\, \$v3534\, \$v2893\, 
               \$v2631\, \$v2669\, \$v3590\, \$v3459\, \$v2695\, \$v2675\, 
               \$v2907\, \$v2898\, \$v2876\, \$v4950\, \$v2811\, \$v2772\, 
               \$v2733\, \$v2808\, \$v2803\, \$v2625\, \$v3422\, \$v2608\, 
               \$v2603\, \$v2567\, \$v2556\, \$v3442\, \$v4994\, \$v2633\, 
               \$v2754\, \$v2602\, \$v2639\, \$v2582\, \$v2829\, \$v2638\, 
               \$v2922\, \$v2792\, \$v5008\, \$v2858\, \$v1527_init\, 
               \$v2743\, \$v1824\, \$v2916\, \$v2779\, \$v3536\, \$v2884\, 
               \$v2817\, \$v2678\, \$v2750\, \$v3517\, \$v2919\, \$v2658\, 
               \$v2891\, \$v2835\, \$v2599\, \$v4974\, \$v2719\, \$v2846\, 
               \$v2805\, \$v2519\, \$v2722\, \$v2865\, \$v2752\, \$v2562\, 
               \$v4924\, \$v2787\, \$v5221\, \$v2874\, \$v2804\, \$v2544\, 
               \$v4944\, \$v2557\, \$v3598\, \$v3518\, rdy1858, \$v2521\, 
               \$v4937\, \$v2756\, \$v3662\, \$v2751\, \$v2744\, \$v3659\, 
               \$v2899\, \$v2825\, \$v2496\, \$v2604\, \$v3605\, \$v2588\, 
               \$v2786\, \$v2522\, \$v3702\, \$v3561\, \$v2877\, \$v2541\, 
               \$v3705\, \$v3602\, \$v2614\, \$v2547\, \$v4991\, \$v2822\, 
               \$v2737\, \$v2640\, \$v4975\, \$v2747\, \$v2553\, \$v1821\, 
               \$v2883\, \$v2610\, \$v3667\, \$v3688\, \$v3607\, \$v2827\, 
               \$v2739\, \$v2713\, \$v2597\, \$v3664\, \$v3472\, \$v2641\, 
               \$v2583\, \$v2525\, \$v2655\, \$v2550\, \$v5017\, \$v2921\, 
               \$v2842\, \$v2710\, \$v3627\, \$v2735\, \$v2689\, \$v2526\, 
               \$v2845\, \$v1815\, \$v2890\, \$v2741\, \$v2612\, \$v3603\, 
               \$v2734\, \$v5029\, \$v2539\, \$v2533\, \$v2757\, \$v2569\, 
               \$v3686\, \$v2511\, \$v2909\, \$v3531\, \$v2702\, \$v2650\, 
               \$v2574\, \$v2502\, \$v4947\, \$v2587\, \$v3624\, \$v2836\, 
               \$v2775\, \$v2624\, \$v2887\, \$v3703\, \$v2694\, \$v2549\, 
               \$v2693\, \$v2634\, \$v2632\, \$v2509\, \$v5306\, \$v2885\, 
               \$v2605\, \$v2558\, \$v2882\, \$v2585\, \$v3613\, \$v3555\
               : value(0 to 0) := (others => '0');
      variable \$711_apply_arg\
               : value(0 to 165) := (others => '0');
      variable \$709_aux_arg\, \$v3479\, \$1050\, \$722_fill_arg\, \$v3468\, 
               \$1052\, \$723_fill_arg\, \$726_w3_arg\
               : value(0 to 79) := (others => '0');
      variable \$719_compbranch_arg\
               : value(0 to 231) := (others => '0');
      variable \$715_binop_compare_arg\
               : value(0 to 153) := (others => '0');
      variable \$5303_v\, \$v5002\, \$5171_v\, \$5482_v\, \$5408\, \$794\, 
               \$1576\, \$5168_v\, \$1616_w\, \$821\, \$5276_v\, 
               compute1859_id, \$5192_v\, \$877_v\, \$1822_v\, \$5499_v\, 
               \$5207_v\, \$5327_v\, \$971_next_env\, \$5544_v\, \$5515_hd\, 
               \$5450\, \$5378_v\, \$1663_hd\, \$1667_hd\, \$5345_v\, 
               \$5383_v\, \$5110_w\, \$5173_v\, \$5363_v\, \$5477_v\, 
               \$5513_v\, \$5316_v\, \$5413\, \$1138\, \$5535_v\, \$5548_v\, 
               \$5137_w\, \$5274_v\, \$5321_v\, \$5325_v\, \$5197_v\, 
               \$5398_v\, \$5263_v\, \$5323_v\, \$5540_v\, \$5202_v\, 
               \$5348_v\, \$5243_v\, \$5336_v\, \$846\, \$5272_v\, \$5306_v\, 
               \$5330_v\, \$5139_hd\, \$5528_v\, \$5295_v\, \$1636\, 
               \$5314_v\, \$788\, \$5403_v\, \$5265_v\, \$5166_v\, \$1104\, 
               \$v4999\, \$1279\, \$5552_v\, \$5351_v\, \$5081_w\, \$5251\, 
               \$5112_hd\, \$5472_v\, \$1235_v\, \$5492_v\, \$5523_v\, 
               \$556_cy\, \$961_f0\, \$5373_v\, \$5542_v\, \$994_next_acc\, 
               \$5550_v\, \$5423\, \$5443\, \$983_v\, \$5360_v\, \$874_v\, 
               \$5467_v\, \$5393_v\, \$5332_v\, \$5436\, \$796_v\, \$v1563\, 
               \$1618_hd\, \$5506_v\, \$5357_v\, \$5418\, \$5311_v\, \$771\, 
               \$1338_v\, \$5429\, \$5530_v\, \$1603\, \$5180_v\, \$1592\, 
               \$5267_v\, \$5388_v\, \$790_v\, \$5334_v\, \$5366_v\, 
               \$5175_v\, \$5318_v\, \$5546_v\, \$1326\, \$5083_hd\, 
               \$5309_v\, \$5354_v\
               : value(0 to 31) := (others => '0');
      variable \$712_offsetclosure_n_result\, \$717_branch_if_result\, 
               \$711_apply_result\, \$716_make_block_n_result\, 
               \$719_compbranch_result\, \$713_binop_int_result\, 
               \$715_binop_compare_result\, \$v8\
               : value(0 to 121) := (others => '0');
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$v3555\); default_zero(\$v3613\); 
          default_zero(\$v2585\); default_zero(\$v2882\); 
          default_zero(\$5354_v\); default_zero(\$v2558\); 
          default_zero(\$v2605\); default_zero(\$v2885\); 
          default_zero(\$v5306\); default_zero(\$v2509\); 
          default_zero(\$v3487\); default_zero(\$v2632\); 
          default_zero(\$v2634\); default_zero(\$v2693\); 
          default_zero(\$5309_v\); default_zero(\$v3611\); 
          default_zero(\$v2549\); default_zero(\$v2694\); 
          default_zero(\$v3703\); default_zero(\$v2887\); 
          default_zero(\$721_w_id\); default_zero(\$v2624\); 
          default_zero(\$v2775\); default_zero(\$v2836\); 
          default_zero(\$5560_sp\); default_zero(\$v3685\); 
          default_zero(\$5083_hd\); default_zero(\$v3624\); 
          default_zero(\$v2587\); default_zero(\$820_sp\); 
          default_zero(\$v4947\); default_zero(\$v2502\); 
          default_zero(\$v2574\); default_zero(\$v2650\); 
          default_zero(\$v2702\); default_zero(\$v3632\); 
          default_zero(\$v3531\); default_zero(\$v3639\); 
          default_zero(\$v2909\); default_zero(\$v2511\); 
          default_zero(\$v3654\); default_zero(\$1326\); 
          default_zero(\$v3686\); default_zero(\$v2569\); 
          default_zero(\$v5300\); default_zero(\$v3600\); 
          default_zero(\$v2757\); default_zero(\$v2533\); 
          default_zero(\$v3646\); default_zero(\$1139_sp\); 
          default_zero(\$v5232\); default_zero(\$v2539\); 
          default_zero(\$v5029\); default_zero(\$v2734\); 
          default_zero(\$v3603\); default_zero(\$v3446\); 
          default_zero(\$5546_v\); default_zero(\$5441_sp\); 
          default_zero(\$v2612\); default_zero(\$v2741\); 
          default_zero(\$v2890\); default_zero(\$5463_sp\); 
          default_zero(\$5318_v\); default_zero(\$v3529\); 
          default_zero(\$v1815\); default_zero(\$v2845\); 
          default_zero(\$v2526\); default_zero(\$v2689\); 
          default_zero(\$v2735\); default_zero(\$v3652\); 
          default_zero(\$5382_sp\); default_zero(\$5175_v\); 
          default_zero(\$v3627\); default_zero(\$5366_v\); 
          default_zero(\$v2710\); default_zero(\$v2842\); 
          default_zero(\$1566\); default_zero(\$5566_sp\); 
          default_zero(\$v2921\); default_zero(\$762_sp\); 
          default_zero(\$v5017\); default_zero(\$713_binop_int_arg\); 
          default_zero(\$5334_v\); default_zero(\$v2550\); 
          default_zero(\$v2655\); default_zero(\$v3551\); 
          default_zero(\$790_v\); default_zero(\$v2525\); 
          default_zero(\$v2583\); default_zero(\$v2641\); 
          default_zero(\$v3472\); default_zero(\$5388_v\); 
          default_zero(\$v3664\); default_zero(\$5267_v\); 
          default_zero(\$v2597\); default_zero(\$v2713\); 
          default_zero(\$v2739\); default_zero(\$v2827\); 
          default_zero(\$v3607\); default_zero(\$v3688\); 
          default_zero(\$717_branch_if_id\); default_zero(\$v3643\); 
          default_zero(\$726_w3_arg\); default_zero(\$1592\); 
          default_zero(\$v3667\); default_zero(\$v2610\); 
          default_zero(\$v2883\); default_zero(\$v1821\); 
          default_zero(\$5180_v\); default_zero(\$v2553\); 
          default_zero(\$v2747\); default_zero(\$1603\); 
          default_zero(\$5530_v\); default_zero(\$v4975\); 
          default_zero(\$v2640\); default_zero(\$903_sp\); 
          default_zero(\$v3640\); default_zero(\$5429\); 
          default_zero(\$v2737\); default_zero(\$v2822\); 
          default_zero(\$1338_v\); default_zero(\$v4991\); 
          default_zero(\$v2547\); default_zero(\$771\); 
          default_zero(\$v2614\); default_zero(\$v3602\); 
          default_zero(\$v3705\); default_zero(\$v2541\); 
          default_zero(\$715_binop_compare_id\); default_zero(\$5377_sp\); 
          default_zero(\$v2877\); default_zero(\$v3561\); 
          default_zero(\$5141\); default_zero(\$v3702\); 
          default_zero(\$v2522\); default_zero(\$v2786\); 
          default_zero(\$819_sp\); default_zero(\$5311_v\); 
          default_zero(\$1581_next\); default_zero(\$v2588\); 
          default_zero(\$894_sp\); default_zero(\$v3605\); 
          default_zero(\$723_fill_arg\); default_zero(\$v2604\); 
          default_zero(\$v2496\); default_zero(\$5563_sp\); 
          default_zero(\$v2825\); default_zero(\$v2899\); 
          default_zero(\$v3659\); default_zero(\$v2744\); 
          default_zero(\$v2751\); default_zero(\$v3662\); 
          default_zero(\$1276_sp\); default_zero(\$v2756\); 
          default_zero(\$v4937\); default_zero(\$v2521\); 
          default_zero(rdy1858); default_zero(\$v3518\); 
          default_zero(\$v3598\); default_zero(\$v2557\); 
          default_zero(\$5418\); default_zero(\$v4944\); 
          default_zero(\$5085\); default_zero(\$5357_v\); 
          default_zero(\$v2544\); default_zero(\$v2804\); 
          default_zero(\$v2874\); default_zero(\$v5221\); 
          default_zero(\$v2787\); default_zero(\$v4924\); 
          default_zero(\$v2562\); default_zero(\$v2752\); 
          default_zero(\$v2865\); default_zero(\$5506_v\); 
          default_zero(\$v2722\); default_zero(\$v2519\); 
          default_zero(\$v2805\); default_zero(\$v2846\); 
          default_zero(\$v2719\); default_zero(\$710_result\); 
          default_zero(\$752_sp\); default_zero(\$v4974\); 
          default_zero(\$v2599\); default_zero(\$v2835\); 
          default_zero(\$v2891\); default_zero(\$v2658\); 
          default_zero(\$v2919\); default_zero(\$v3517\); 
          default_zero(\$v2750\); default_zero(\$v3700\); 
          default_zero(\$v3622\); default_zero(\$v2678\); 
          default_zero(\$v2817\); default_zero(\$v2884\); 
          default_zero(\$v3536\); default_zero(\$1275_sp\); 
          default_zero(\$v2779\); default_zero(\$v2916\); 
          default_zero(\$v1824\); default_zero(\$v2743\); 
          default_zero(\$v1527_init\); default_zero(\$v3683\); 
          default_zero(\$v2858\); default_zero(\$875_sp\); 
          default_zero(\$1618_hd\); default_zero(\$721_w_arg\); 
          default_zero(\$v1563\); default_zero(\$v5008\); 
          default_zero(\$v2792\); default_zero(\$v2922\); 
          default_zero(\$v2638\); default_zero(\$v2829\); 
          default_zero(\$v2582\); default_zero(\$796_v\); 
          default_zero(\$v2639\); default_zero(\$5436\); 
          default_zero(\$v2602\); default_zero(\$v2754\); 
          default_zero(\$970_sp\); default_zero(\$709_aux_id\); 
          default_zero(\$v2633\); default_zero(\$v3690\); 
          default_zero(\$v4994\); default_zero(\$1277_sp\); 
          default_zero(\$v3442\); default_zero(\$v2556\); 
          default_zero(\$724_w0_id\); default_zero(\$713_binop_int_id\); 
          default_zero(\$744_argument1\); default_zero(\$5332_v\); 
          default_zero(\$717_branch_if_arg\); default_zero(\$v2567\); 
          default_zero(\$5393_v\); default_zero(\$724_w0_result\); 
          default_zero(\$715_binop_compare_arg\); default_zero(\$v2603\); 
          default_zero(\$v2608\); default_zero(\$5467_v\); 
          default_zero(\$902_sp\); default_zero(\$718_loop_push_id\); 
          default_zero(\$v1820\); default_zero(\$5114\); 
          default_zero(\$v3422\); default_zero(\$v2625\); 
          default_zero(\$v2803\); default_zero(\$v3645\); 
          default_zero(\$1565_next\); default_zero(\$v2808\); 
          default_zero(\$v8\); default_zero(\$v2733\); 
          default_zero(\$v2772\); default_zero(\$v2811\); 
          default_zero(\$874_v\); default_zero(\$714_compare_arg\); 
          default_zero(\$v4950\); default_zero(\$v2876\); 
          default_zero(\$v2898\); default_zero(\$747\); 
          default_zero(\$v2907\); default_zero(\$v2675\); 
          default_zero(\$v2695\); default_zero(\$v3459\); 
          default_zero(\$v3590\); default_zero(\$v2669\); 
          default_zero(\$1055\); default_zero(\$5360_v\); 
          default_zero(\$v3486\); default_zero(\$v2631\); 
          default_zero(\$v2893\); default_zero(\$v3534\); 
          default_zero(\$v3669\); default_zero(\$v2864\); 
          default_zero(\$v2611\); default_zero(\$v2690\); 
          default_zero(\$936_sp\); default_zero(\$983_v\); 
          default_zero(\$723_fill_result\); default_zero(\$v2584\); 
          default_zero(\$v3542\); default_zero(\$719_compbranch_arg\); 
          default_zero(\$v3419\); default_zero(\$1218_res\); 
          default_zero(\$v2715\); default_zero(\$v3647\); 
          default_zero(\$706_loop_arg\); default_zero(rdy4919); 
          default_zero(\$v3608\); default_zero(\$v2673\); 
          default_zero(\$v5304\); default_zero(\$v3692\); 
          default_zero(\$v3597\); default_zero(\$v4965\); 
          default_zero(\$v2590\); default_zero(\$1284_sp\); 
          default_zero(\$v3505\); default_zero(\$v5297\); 
          default_zero(\$v3591\); default_zero(\$v1822\); 
          default_zero(\$5443\); default_zero(\$v2527\); 
          default_zero(\$v2560\); default_zero(\$720_w_id\); 
          default_zero(\$711_apply_id\); default_zero(\$5423\); 
          default_zero(\$v2671\); default_zero(\$v2793\); 
          default_zero(\$v3657\); default_zero(\$v3419_init\); 
          default_zero(\$v3594\); default_zero(\$714_compare_id\); 
          default_zero(\$v2749\); default_zero(\$5387_sp\); 
          default_zero(\$1052\); default_zero(\$v3673\); 
          default_zero(\$v3650\); default_zero(\$v2813\); 
          default_zero(\$v2839\); default_zero(\$5550_v\); 
          default_zero(\$v2742\); default_zero(\$v2918\); 
          default_zero(\$v3704\); default_zero(\$715_binop_compare_result\); 
          default_zero(\$v2619\); default_zero(\$v2852\); 
          default_zero(\$994_next_acc\); default_zero(\$v2665\); 
          default_zero(\$v2855\); default_zero(\$5542_v\); 
          default_zero(\$710_arg\); default_zero(\$v1549\); 
          default_zero(\$v2753\); default_zero(\$1332_sp\); 
          default_zero(\$v2662\); default_zero(\$v2902\); 
          default_zero(\$v3564\); default_zero(\$v3644\); 
          default_zero(\$v3681\); default_zero(\$5557_sp\); 
          default_zero(\$923_sp\); default_zero(\$5373_v\); 
          default_zero(\$v2724\); default_zero(\$v2915\); 
          default_zero(\$5427_sp\); default_zero(\$912_sp\); 
          default_zero(\$v3506\); default_zero(\$v2629\); 
          default_zero(\$v2648\); default_zero(\$v2616\); 
          default_zero(\$v2736\); default_zero(\$v3696\); 
          default_zero(\$961_f0\); default_zero(\$v2821\); 
          default_zero(\$v3460\); default_zero(\$v5294\); 
          default_zero(\$v3593\); default_zero(\$v2672\); 
          default_zero(\$v3668\); default_zero(\$v2925\); 
          default_zero(\$v2512\); default_zero(\$v4984\); 
          default_zero(\$5372_sp\); default_zero(\$v2552\); 
          default_zero(\$v2618\); default_zero(\$v2911\); 
          default_zero(\$556_cy\); default_zero(\$5523_v\); 
          default_zero(\$5492_v\); default_zero(\$v2738\); 
          default_zero(\$v3623\); default_zero(\$712_offsetclosure_n_arg\); 
          default_zero(\$v2685\); default_zero(\$v2859\); 
          default_zero(\$v3552\); default_zero(\$1235_v\); 
          default_zero(\$5472_v\); default_zero(\$v2555\); 
          default_zero(\$725_w1_id\); default_zero(\$5112_hd\); 
          default_zero(\$v3447\); default_zero(\$5251\); 
          default_zero(\$v2778\); default_zero(\$v2802\); 
          default_zero(\$764_sp\); default_zero(\$v3615\); 
          default_zero(\$v3576\); default_zero(\$v2623\); 
          default_zero(\$v2637\); default_zero(\$721_w_result\); 
          default_zero(\$v2771\); default_zero(\$v2853\); 
          default_zero(\$v2888\); default_zero(\$v3628\); 
          default_zero(\$5081_w\); default_zero(\$v2621\); 
          default_zero(\$5351_v\); default_zero(\$v3675\); 
          default_zero(\$v2682\); default_zero(\$v3638\); 
          default_zero(\$v4997\); default_zero(\$v2819\); 
          default_zero(\$v3589\); default_zero(\$v2663\); 
          default_zero(\$v2814\); default_zero(\$726_w3_id\); 
          default_zero(\$v3691\); default_zero(\$v2716\); 
          default_zero(\$1620\); default_zero(\$5552_v\); 
          default_zero(\$v2528\); default_zero(\$v2666\); 
          default_zero(\$v2703\); default_zero(\$v2559\); 
          default_zero(\$v2755\); default_zero(\$v3618\); 
          default_zero(\$5434_sp\); default_zero(\$v3530\); 
          default_zero(\$v2929\); default_zero(\$v2576\); 
          default_zero(\$v3658\); default_zero(\$v2850\); 
          default_zero(\$v2863\); default_zero(\$1279\); 
          default_zero(\$v2816\); default_zero(\$708_loop_id\); 
          default_zero(\$v2654\); default_zero(\$v1545_init\); 
          default_zero(\$v2613\); default_zero(\$v2758\); 
          default_zero(\$713_binop_int_result\); 
          default_zero(\$719_compbranch_result\); default_zero(\$v2677\); 
          default_zero(\$v2880\); default_zero(\$v3533\); 
          default_zero(\$v2532\); default_zero(\$v2698\); 
          default_zero(\$v2886\); default_zero(\$v4999\); 
          default_zero(\$v2770\); default_zero(\$1104\); 
          default_zero(\$v2537\); default_zero(\$5166_v\); 
          default_zero(\$5265_v\); default_zero(\$v2538\); 
          default_zero(\$v3612\); default_zero(\$v3468\); 
          default_zero(\$5403_v\); default_zero(\$v2878\); 
          default_zero(\$v2881\); default_zero(\$v3572\); 
          default_zero(\$788\); default_zero(\$5314_v\); 
          default_zero(\$724_w0_arg\); default_zero(\$v2571\); 
          default_zero(\$v2647\); default_zero(\$v2668\); 
          default_zero(\$1636\); default_zero(\$v3596\); 
          default_zero(\$v2529\); default_zero(\$v2810\); 
          default_zero(\$v3616\); default_zero(\$v3697\); 
          default_zero(\$v2840\); default_zero(\$v5012\); 
          default_zero(\$v2535\); default_zero(\$v2595\); 
          default_zero(\$v2777\); default_zero(\$v3570\); 
          default_zero(\$708_loop_arg\); default_zero(\$v2828\); 
          default_zero(\$901_sp\); default_zero(\$v3620\); 
          default_zero(\$778_sp\); default_zero(\$v3655\); 
          default_zero(\$v2507\); default_zero(\$v2615\); 
          default_zero(\$v1825\); default_zero(\$v5194\); 
          default_zero(\$v2659\); default_zero(\$v2717\); 
          default_zero(\$v2851\); default_zero(\$v2871\); 
          default_zero(\$888_idx\); default_zero(\$v2667\); 
          default_zero(\$5295_v\); default_zero(\$5528_v\); 
          default_zero(\$5139_hd\); default_zero(\$5330_v\); 
          default_zero(\$5306_v\); default_zero(\$v2657\); 
          default_zero(\$v2906\); default_zero(\$745_argument2\); 
          default_zero(\$v3699\); default_zero(\$v5037\); 
          default_zero(\$v1810\); default_zero(\$v2628\); 
          default_zero(\$v2718\); default_zero(\$5272_v\); 
          default_zero(\$1305_sp\); default_zero(\$846\); 
          default_zero(\$v2499\); default_zero(\$v2506\); 
          default_zero(\$v2561\); default_zero(\$v2732\); 
          default_zero(\$v3689\); default_zero(\$v3701\); 
          default_zero(\$709_aux_result\); default_zero(\$v2600\); 
          default_zero(\$v3478\); default_zero(\$v2745\); 
          default_zero(\$v2784\); default_zero(\$v2551\); 
          default_zero(\$v2593\); default_zero(\$v2785\); 
          default_zero(\$v2504\); default_zero(\$v2606\); 
          default_zero(\$v3573\); default_zero(\$5336_v\); 
          default_zero(\$v2913\); default_zero(\$763_sp\); 
          default_zero(\$v3619\); default_zero(\$v2856\); 
          default_zero(\$v2903\); default_zero(\$v2746\); 
          default_zero(\$v2815\); default_zero(\$v2643\); 
          default_zero(\$v2661\); default_zero(\$v3547\); 
          default_zero(\$v2642\); default_zero(\$v3535\); 
          default_zero(\$v3671\); default_zero(\$v3663\); 
          default_zero(\$707_copy_root_in_ram_result\); 
          default_zero(\$v2708\); default_zero(\$5243_v\); 
          default_zero(\$v2572\); default_zero(\$v2830\); 
          default_zero(\$v1563_init\); default_zero(\$v3672\); 
          default_zero(\$v3516\); default_zero(\$v2759\); 
          default_zero(\$v3614\); default_zero(\$5348_v\); 
          default_zero(\$v2794\); default_zero(\$5402_sp\); 
          default_zero(\$v2709\); default_zero(\$1312_sp\); 
          default_zero(\$5202_v\); default_zero(\$722_fill_arg\); 
          default_zero(\$v2826\); default_zero(\$v2620\); 
          default_zero(\$v2857\); default_zero(\$712_offsetclosure_n_id\); 
          default_zero(\$5540_v\); default_zero(\$v2924\); 
          default_zero(\$v2645\); default_zero(\$814_sp\); 
          default_zero(\$v5033\); default_zero(\$v2807\); 
          default_zero(\$v2843\); default_zero(\$1180_sp\); 
          default_zero(\$v2797\); default_zero(\$708_loop_result\); 
          default_zero(\$v2849\); default_zero(\$1530\); 
          default_zero(\$v2799\); default_zero(\$v2895\); 
          default_zero(\$v3666\); default_zero(\$v2591\); 
          default_zero(\$1038_sp\); default_zero(\$v2847\); 
          default_zero(\$v5311\); default_zero(\$976\); 
          default_zero(\$v2510\); default_zero(\$v3682\); 
          default_zero(\$v2767\); default_zero(\$v3625\); 
          default_zero(\$v5288\); default_zero(\$v2622\); 
          default_zero(\$v2841\); default_zero(\$v2892\); 
          default_zero(\$707_copy_root_in_ram_id\); default_zero(\$v2831\); 
          default_zero(\$v2917\); default_zero(\$v2577\); 
          default_zero(\$v5228\); default_zero(\$v2554\); 
          default_zero(\$v2832\); default_zero(\$v2896\); 
          default_zero(\$v2697\); default_zero(\$v2518\); 
          default_zero(\$547_o\); default_zero(\$v2601\); 
          default_zero(\$v2598\); default_zero(\$v3633\); 
          default_zero(\$v2575\); default_zero(\$5323_v\); 
          default_zero(\$1196_res\); default_zero(\$v2596\); 
          default_zero(\$v2644\); default_zero(\$v2536\); 
          default_zero(\$v2681\); default_zero(\$v3601\); 
          default_zero(\$v3637\); default_zero(rdy2975); 
          default_zero(\$722_fill_id\); default_zero(\$5263_v\); 
          default_zero(\$v1557\); default_zero(\$v2586\); 
          default_zero(\$785_sp\); default_zero(\$v2867\); 
          default_zero(\$v1545\); default_zero(\$v2570\); 
          default_zero(\$716_make_block_n_result\); default_zero(\$v2515\); 
          default_zero(result2974); default_zero(\$v5041\); 
          default_zero(\$v3528\); default_zero(\$v2692\); 
          default_zero(\$v2872\); default_zero(\$v3634\); 
          default_zero(\$v2727\); default_zero(\$v4962\); 
          default_zero(\$v3545\); default_zero(\$879_sp\); 
          default_zero(\$718_loop_push_arg\); default_zero(\$v2676\); 
          default_zero(\$710_id\); default_zero(\$v3604\); 
          default_zero(\$5398_v\); default_zero(\$720_w_arg\); 
          default_zero(\$v2683\); default_zero(\$v2711\); 
          default_zero(\$v2763\); default_zero(\$726_w3_result\); 
          default_zero(\$716_make_block_n_arg\); default_zero(\$v3443\); 
          default_zero(\$5197_v\); default_zero(\$5325_v\); 
          default_zero(\$v2927\); default_zero(\$v495\); 
          default_zero(\$v2568\); default_zero(\$v2578\); 
          default_zero(\$v2908\); default_zero(\$v3558\); 
          default_zero(\$v2720\); default_zero(\$v2721\); 
          default_zero(\$v3503\); default_zero(\$1243_sp\); 
          default_zero(\$v2609\); default_zero(\$5321_v\); 
          default_zero(\$v4988\); default_zero(\$5274_v\); 
          default_zero(\$v2705\); default_zero(\$v2861\); 
          default_zero(\$v4982\); default_zero(\$711_apply_arg\); 
          default_zero(\$v1860\); default_zero(\$v3444\); 
          default_zero(\$718_loop_push_result\); default_zero(\$v3504\); 
          default_zero(\$v2626\); default_zero(\$v5246\); 
          default_zero(\$v2565\); default_zero(\$v2740\); 
          default_zero(\$5397_sp\); default_zero(\$1568_next\); 
          default_zero(\$v3563\); default_zero(\$v3649\); 
          default_zero(\$v3629\); default_zero(\$v2848\); 
          default_zero(\$v2860\); default_zero(\$720_w_result\); 
          default_zero(\$v3458\); default_zero(\$v2548\); 
          default_zero(\$v2563\); default_zero(\$v2686\); 
          default_zero(\$v2765\); default_zero(\$v1814\); 
          default_zero(\$5137_w\); default_zero(\$v5048\); 
          default_zero(\$v4998\); default_zero(\$5548_v\); 
          default_zero(\$v2862\); default_zero(\$5535_v\); 
          default_zero(\$v2930\); default_zero(\$v2530\); 
          default_zero(\$v2823\); default_zero(\$v3676\); 
          default_zero(\$v2869\); default_zero(\$1138\); 
          default_zero(\$v3684\); default_zero(\$v5308\); 
          default_zero(\$v2795\); default_zero(\$v2889\); 
          default_zero(\$v2723\); default_zero(\$v2517\); 
          default_zero(\$v5238\); default_zero(\$v2904\); 
          default_zero(\$5461_sp\); default_zero(\$5413\); 
          default_zero(\$v2905\); default_zero(\$v3631\); 
          default_zero(\$v2684\); default_zero(\$v2696\); 
          default_zero(\$v5025\); default_zero(\$1278_sp\); 
          default_zero(\$v2824\); default_zero(\$v2834\); 
          default_zero(\$v2514\); default_zero(\$723_fill_id\); 
          default_zero(\$v2531\); default_zero(\$v2920\); 
          default_zero(\$v2573\); default_zero(\$v3519\); 
          default_zero(\$v1823\); default_zero(\$1288_sp\); 
          default_zero(\$5316_v\); default_zero(\$v3665\); 
          default_zero(\$v1549_init\); default_zero(\$v3670\); 
          default_zero(\$v2579\); default_zero(\$v3549\); 
          default_zero(\$1179_sp\); default_zero(\$883_ofs\); 
          default_zero(\$v4980\); default_zero(\$v2932\); 
          default_zero(\$v2806\); default_zero(\$5513_v\); 
          default_zero(\$5392_sp\); default_zero(\$v2664\); 
          default_zero(\$v3595\); default_zero(\$v2687\); 
          default_zero(\$v2701\); default_zero(\$v2766\); 
          default_zero(\$v2729\); default_zero(\$v3698\); 
          default_zero(\$v2636\); default_zero(\$v2594\); 
          default_zero(\$v2679\); default_zero(\$v2699\); 
          default_zero(\$v2790\); default_zero(\$5477_v\); 
          default_zero(\$v2926\); default_zero(\$v2497\); 
          default_zero(\$5448_sp\); default_zero(\$v2789\); 
          default_zero(\$v2798\); default_zero(\$v3592\); 
          default_zero(\$v4931\); default_zero(\$792_sp\); 
          default_zero(\$v5291\); default_zero(\$v4953\); 
          default_zero(\$1101\); default_zero(\$v3427\); 
          default_zero(\$v3653\); default_zero(\$707_copy_root_in_ram_arg\); 
          default_zero(\$v2589\); default_zero(\$v2707\); 
          default_zero(\$711_apply_result\); default_zero(\$5363_v\); 
          default_zero(\$v2674\); default_zero(\$v2760\); 
          default_zero(\$v2566\); default_zero(\$5173_v\); 
          default_zero(\$v2776\); default_zero(\$v3642\); 
          default_zero(\$v2543\); default_zero(\$v2773\); 
          default_zero(\$5110_w\); default_zero(\$v3626\); 
          default_zero(\$v2635\); default_zero(\$1152_arg\); 
          default_zero(\$v2870\); default_zero(\$5383_v\); 
          default_zero(\$v1808\); default_zero(\$v2649\); 
          default_zero(\$v2706\); default_zero(\$5345_v\); 
          default_zero(\$v3661\); default_zero(\$v2796\); 
          default_zero(\$v3610\); default_zero(\$v5046\); 
          default_zero(\$v2680\); default_zero(\$725_w1_arg\); 
          default_zero(\$v2910\); default_zero(\$v3617\); 
          default_zero(\$893_sp\); default_zero(\$719_compbranch_id\); 
          default_zero(\$1567_next\); default_zero(\$v1557_init\); 
          default_zero(\$v2728\); default_zero(\$v2546\); 
          default_zero(\$v2894\); default_zero(\$v3415\); 
          default_zero(\$v3550\); default_zero(\$1667_hd\); 
          default_zero(\$v2688\); default_zero(\$v2838\); 
          default_zero(\$859_sp\); default_zero(\$706_loop_result\); 
          default_zero(\$1663_hd\); default_zero(\$706_loop_id\); 
          default_zero(\$v5307\); default_zero(\$v2933\); 
          default_zero(\$v2901\); default_zero(\$v2523\); 
          default_zero(\$v2780\); default_zero(\$5378_v\); 
          default_zero(\$v2524\); default_zero(\$v2700\); 
          default_zero(\$5450\); default_zero(\$v2833\); 
          default_zero(\$v2900\); default_zero(\$v2542\); 
          default_zero(\$v2714\); default_zero(\$1285_sp\); 
          default_zero(\$1297_sp\); default_zero(\$717_branch_if_result\); 
          default_zero(\$v2879\); default_zero(\$v3457\); 
          default_zero(\$5515_hd\); default_zero(\$1050\); 
          default_zero(\$v2503\); default_zero(\$5544_v\); 
          default_zero(\$v3695\); default_zero(\$v2725\); 
          default_zero(\$v2508\); default_zero(\$v2704\); 
          default_zero(\$v3477\); default_zero(\$v2923\); 
          default_zero(\$v2564\); default_zero(\$v2914\); 
          default_zero(\$v3660\); default_zero(\$971_next_env\); 
          default_zero(\$v2691\); default_zero(\$5327_v\); 
          default_zero(\$v2801\); default_zero(\$5207_v\); 
          default_zero(\$v3636\); 
          default_zero(\$712_offsetclosure_n_result\); 
          default_zero(\$5499_v\); default_zero(\$v2800\); 
          default_zero(\$1822_v\); default_zero(\$v1556_init\); 
          default_zero(\$v2837\); default_zero(\$v2500\); 
          default_zero(\$v5256\); default_zero(\$877_v\); 
          default_zero(\$v2513\); default_zero(\$5370_sp\); 
          default_zero(\$v2761\); default_zero(\$v2844\); 
          default_zero(\$v2897\); default_zero(\$v2912\); 
          default_zero(\$v3674\); default_zero(\$v2818\); 
          default_zero(\$5192_v\); default_zero(\$1127_b\); 
          default_zero(\$v2581\); default_zero(\$v2656\); 
          default_zero(\$v2873\); default_zero(result1857); 
          default_zero(compute1859_id); default_zero(\$v3606\); 
          default_zero(\$v3694\); default_zero(\$v2782\); 
          default_zero(\$v2866\); default_zero(\$v2545\); 
          default_zero(\$v3559\); default_zero(\$v5303\); 
          default_zero(\$v2931\); default_zero(\$v2712\); 
          default_zero(\$v14\); default_zero(\$v3599\); 
          default_zero(\$v2670\); default_zero(\$722_fill_result\); 
          default_zero(\$v2627\); default_zero(\$v3693\); 
          default_zero(\$v4971\); default_zero(\$v3441\); 
          default_zero(\$v232\); default_zero(\$v2630\); 
          default_zero(\$v3575\); default_zero(\$v3416\); 
          default_zero(\$5276_v\); default_zero(\$v2540\); 
          default_zero(\$v3479\); default_zero(\$v5310\); 
          default_zero(\$951_sp\); default_zero(\$v2726\); 
          default_zero(\$821\); default_zero(\$v2607\); 
          default_zero(\$725_w1_result\); default_zero(\$v2646\); 
          default_zero(\$v2651\); default_zero(\$v3651\); 
          default_zero(\$967\); default_zero(\$803_sp\); 
          default_zero(\$v2730\); default_zero(\$1616_w\); 
          default_zero(\$v2788\); default_zero(\$v2660\); 
          default_zero(\$5168_v\); default_zero(\$740\); 
          default_zero(\$714_compare_result\); default_zero(\$v2653\); 
          default_zero(\$v2781\); default_zero(\$v2875\); 
          default_zero(\$885\); default_zero(result4918); 
          default_zero(\$v1527\); default_zero(\$v1818\); 
          default_zero(\$v5203\); default_zero(\$v3687\); 
          default_zero(\$1579\); default_zero(\$v3609\); 
          default_zero(\$548_rdy\); default_zero(\$v2520\); 
          default_zero(\$v2731\); default_zero(\$v3567\); 
          default_zero(\$v2783\); default_zero(\$v3548\); 
          default_zero(\$v5274\); default_zero(\$v2505\); 
          default_zero(\$v2617\); default_zero(\$v2768\); 
          default_zero(\$v2762\); default_zero(\$v2854\); 
          default_zero(\$1576\); default_zero(\$975_sp\); 
          default_zero(\$716_make_block_n_id\); default_zero(\$v2812\); 
          default_zero(\$v3417\); default_zero(\$v1809\); 
          default_zero(\$v2764\); default_zero(\$v3532\); 
          default_zero(\$v2774\); default_zero(\$v2809\); 
          default_zero(\$v5014\); default_zero(\$794\); 
          default_zero(\$5408\); default_zero(\$v2748\); 
          default_zero(\$v3566\); default_zero(\$v4976\); 
          default_zero(\$v2791\); default_zero(\$5482_v\); 
          default_zero(\$v1556\); default_zero(\$746_argument3\); 
          default_zero(\$709_aux_arg\); default_zero(\$v2592\); 
          default_zero(\$v2580\); default_zero(\$v3569\); 
          default_zero(\$5171_v\); default_zero(\$v2868\); 
          default_zero(\$v4934\); default_zero(\$v5002\); 
          default_zero(\$v2652\); default_zero(\$v3428\); 
          default_zero(\$v2516\); default_zero(\$5459_sp\); 
          default_zero(\$v2928\); default_zero(\$v2534\); 
          default_zero(\$v2820\); default_zero(\$v2769\); 
          default_zero(\$5303_v\); default_zero(\$v5021\); 
          default_zero(\$v2498\); default_zero(\$v2501\); 
          default_zero(\$v5309\); 
          rdy <= "1";
          rdy1858 := "0";
          state <= compute1859;
          state_var5313 <= compute2976;
          state_var5312 <= compute4920;
          
        else if run = '1' then
          case state is
          when compute1859 =>
            rdy1858 := eclat_false;
            \$v5311\ := eclat_not(\$v1563_init\);
            if \$v5311\(0) = '1' then
              \$v1563\ := X"0000000" & X"0";
              \$v1563_init\ := eclat_true;
            end if;
            \$v1563\ := eclat_if(eclat_false & X"0000000" & X"0" & eclat_add(\$v1563\ & X"0000000" & X"1"));
            \$v1825\ := eclat_unit;
            \$556_cy\ := \$v1563\;
            \$v5310\ := eclat_not(\$v1527_init\);
            if \$v5310\(0) = '1' then
              \$v1527\ := eclat_false & eclat_false & eclat_false & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_false;
              \$v1527_init\ := eclat_true;
            end if;
            \$v5309\ := eclat_not(""&\$v1527\(2));
            if \$v5309\(0) = '1' then
              \$v3415\ := eclat_not(\$v1557_init\);
              if \$v3415\(0) = '1' then
                \$v1557\ := eclat_unit & eclat_false;
                \$v1557_init\ := eclat_true;
              end if;
              case state_var5313 is
              when pause_setI2977 =>
                \$code_write_request\ <= '0';
                \$v2919\ := eclat_unit;
                \$v14\ := eclat_unit;
                \$v1557\ := \$v14\ & eclat_true;
                result2974 := eclat_unit;
                rdy2975 := eclat_true;
                state_var5313 <= compute2976;
              when pause_setI2978 =>
                \$code_write_request\ <= '0';
                \$v2918\ := eclat_unit;
                \$code_ptr_write\ <= 421;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"8f";
                state_var5313 <= pause_setI2977;
              when pause_setI2979 =>
                \$code_write_request\ <= '0';
                \$v2917\ := eclat_unit;
                \$code_ptr_write\ <= 420;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"5";
                state_var5313 <= pause_setI2978;
              when pause_setI2980 =>
                \$code_write_request\ <= '0';
                \$v2916\ := eclat_unit;
                \$code_ptr_write\ <= 419;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"13";
                state_var5313 <= pause_setI2979;
              when pause_setI2981 =>
                \$code_write_request\ <= '0';
                \$v2915\ := eclat_unit;
                \$code_ptr_write\ <= 418;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI2980;
              when pause_setI2982 =>
                \$code_write_request\ <= '0';
                \$v2914\ := eclat_unit;
                \$code_ptr_write\ <= 417;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"13";
                state_var5313 <= pause_setI2981;
              when pause_setI2983 =>
                \$code_write_request\ <= '0';
                \$v2913\ := eclat_unit;
                \$code_ptr_write\ <= 416;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"e");
                state_var5313 <= pause_setI2982;
              when pause_setI2984 =>
                \$code_write_request\ <= '0';
                \$v2912\ := eclat_unit;
                \$code_ptr_write\ <= 415;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"55";
                state_var5313 <= pause_setI2983;
              when pause_setI2985 =>
                \$code_write_request\ <= '0';
                \$v2911\ := eclat_unit;
                \$code_ptr_write\ <= 414;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7a";
                state_var5313 <= pause_setI2984;
              when pause_setI2986 =>
                \$code_write_request\ <= '0';
                \$v2910\ := eclat_unit;
                \$code_ptr_write\ <= 413;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI2985;
              when pause_setI2987 =>
                \$code_write_request\ <= '0';
                \$v2909\ := eclat_unit;
                \$code_ptr_write\ <= 412;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI2986;
              when pause_setI2988 =>
                \$code_write_request\ <= '0';
                \$v2908\ := eclat_unit;
                \$code_ptr_write\ <= 411;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"14";
                state_var5313 <= pause_setI2987;
              when pause_setI2989 =>
                \$code_write_request\ <= '0';
                \$v2907\ := eclat_unit;
                \$code_ptr_write\ <= 410;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI2988;
              when pause_setI2990 =>
                \$code_write_request\ <= '0';
                \$v2906\ := eclat_unit;
                \$code_ptr_write\ <= 409;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7f";
                state_var5313 <= pause_setI2989;
              when pause_setI2991 =>
                \$code_write_request\ <= '0';
                \$v2905\ := eclat_unit;
                \$code_ptr_write\ <= 408;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"9";
                state_var5313 <= pause_setI2990;
              when pause_setI2992 =>
                \$code_write_request\ <= '0';
                \$v2904\ := eclat_unit;
                \$code_ptr_write\ <= 407;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI2991;
              when pause_setI2993 =>
                \$code_write_request\ <= '0';
                \$v2903\ := eclat_unit;
                \$code_ptr_write\ <= 406;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI2992;
              when pause_setI2994 =>
                \$code_write_request\ <= '0';
                \$v2902\ := eclat_unit;
                \$code_ptr_write\ <= 405;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI2993;
              when pause_setI2995 =>
                \$code_write_request\ <= '0';
                \$v2901\ := eclat_unit;
                \$code_ptr_write\ <= 404;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"7";
                state_var5313 <= pause_setI2994;
              when pause_setI2996 =>
                \$code_write_request\ <= '0';
                \$v2900\ := eclat_unit;
                \$code_ptr_write\ <= 403;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"67";
                state_var5313 <= pause_setI2995;
              when pause_setI2997 =>
                \$code_write_request\ <= '0';
                \$v2899\ := eclat_unit;
                \$code_ptr_write\ <= 402;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"5c";
                state_var5313 <= pause_setI2996;
              when pause_setI2998 =>
                \$code_write_request\ <= '0';
                \$v2898\ := eclat_unit;
                \$code_ptr_write\ <= 401;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"10";
                state_var5313 <= pause_setI2997;
              when pause_setI2999 =>
                \$code_write_request\ <= '0';
                \$v2897\ := eclat_unit;
                \$code_ptr_write\ <= 400;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"55";
                state_var5313 <= pause_setI2998;
              when pause_setI3000 =>
                \$code_write_request\ <= '0';
                \$v2896\ := eclat_unit;
                \$code_ptr_write\ <= 399;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7d";
                state_var5313 <= pause_setI2999;
              when pause_setI3001 =>
                \$code_write_request\ <= '0';
                \$v2895\ := eclat_unit;
                \$code_ptr_write\ <= 398;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3000;
              when pause_setI3002 =>
                \$code_write_request\ <= '0';
                \$v2894\ := eclat_unit;
                \$code_ptr_write\ <= 397;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"9";
                state_var5313 <= pause_setI3001;
              when pause_setI3003 =>
                \$code_write_request\ <= '0';
                \$v2893\ := eclat_unit;
                \$code_ptr_write\ <= 396;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"69";
                state_var5313 <= pause_setI3002;
              when pause_setI3004 =>
                \$code_write_request\ <= '0';
                \$v2892\ := eclat_unit;
                \$code_ptr_write\ <= 395;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"69";
                state_var5313 <= pause_setI3003;
              when pause_setI3005 =>
                \$code_write_request\ <= '0';
                \$v2891\ := eclat_unit;
                \$code_ptr_write\ <= 394;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"fb");
                state_var5313 <= pause_setI3004;
              when pause_setI3006 =>
                \$code_write_request\ <= '0';
                \$v2890\ := eclat_unit;
                \$code_ptr_write\ <= 393;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3005;
              when pause_setI3007 =>
                \$code_write_request\ <= '0';
                \$v2889\ := eclat_unit;
                \$code_ptr_write\ <= 392;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3006;
              when pause_setI3008 =>
                \$code_write_request\ <= '0';
                \$v2888\ := eclat_unit;
                \$code_ptr_write\ <= 391;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"13";
                state_var5313 <= pause_setI3007;
              when pause_setI3009 =>
                \$code_write_request\ <= '0';
                \$v2887\ := eclat_unit;
                \$code_ptr_write\ <= 390;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3008;
              when pause_setI3010 =>
                \$code_write_request\ <= '0';
                \$v2886\ := eclat_unit;
                \$code_ptr_write\ <= 389;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"c6");
                state_var5313 <= pause_setI3009;
              when pause_setI3011 =>
                \$code_write_request\ <= '0';
                \$v2885\ := eclat_unit;
                \$code_ptr_write\ <= 388;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3010;
              when pause_setI3012 =>
                \$code_write_request\ <= '0';
                \$v2884\ := eclat_unit;
                \$code_ptr_write\ <= 387;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3011;
              when pause_setI3013 =>
                \$code_write_request\ <= '0';
                \$v2883\ := eclat_unit;
                \$code_ptr_write\ <= 386;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"f";
                state_var5313 <= pause_setI3012;
              when pause_setI3014 =>
                \$code_write_request\ <= '0';
                \$v2882\ := eclat_unit;
                \$code_ptr_write\ <= 385;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3013;
              when pause_setI3015 =>
                \$code_write_request\ <= '0';
                \$v2881\ := eclat_unit;
                \$code_ptr_write\ <= 384;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"9b");
                state_var5313 <= pause_setI3014;
              when pause_setI3016 =>
                \$code_write_request\ <= '0';
                \$v2880\ := eclat_unit;
                \$code_ptr_write\ <= 383;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3015;
              when pause_setI3017 =>
                \$code_write_request\ <= '0';
                \$v2879\ := eclat_unit;
                \$code_ptr_write\ <= 382;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3016;
              when pause_setI3018 =>
                \$code_write_request\ <= '0';
                \$v2878\ := eclat_unit;
                \$code_ptr_write\ <= 381;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"e";
                state_var5313 <= pause_setI3017;
              when pause_setI3019 =>
                \$code_write_request\ <= '0';
                \$v2877\ := eclat_unit;
                \$code_ptr_write\ <= 380;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3018;
              when pause_setI3020 =>
                \$code_write_request\ <= '0';
                \$v2876\ := eclat_unit;
                \$code_ptr_write\ <= 379;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3019;
              when pause_setI3021 =>
                \$code_write_request\ <= '0';
                \$v2875\ := eclat_unit;
                \$code_ptr_write\ <= 378;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"e";
                state_var5313 <= pause_setI3020;
              when pause_setI3022 =>
                \$code_write_request\ <= '0';
                \$v2874\ := eclat_unit;
                \$code_ptr_write\ <= 377;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"64";
                state_var5313 <= pause_setI3021;
              when pause_setI3023 =>
                \$code_write_request\ <= '0';
                \$v2873\ := eclat_unit;
                \$code_ptr_write\ <= 376;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"10";
                state_var5313 <= pause_setI3022;
              when pause_setI3024 =>
                \$code_write_request\ <= '0';
                \$v2872\ := eclat_unit;
                \$code_ptr_write\ <= 375;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3023;
              when pause_setI3025 =>
                \$code_write_request\ <= '0';
                \$v2871\ := eclat_unit;
                \$code_ptr_write\ <= 374;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"5b");
                state_var5313 <= pause_setI3024;
              when pause_setI3026 =>
                \$code_write_request\ <= '0';
                \$v2870\ := eclat_unit;
                \$code_ptr_write\ <= 373;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3025;
              when pause_setI3027 =>
                \$code_write_request\ <= '0';
                \$v2869\ := eclat_unit;
                \$code_ptr_write\ <= 372;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3026;
              when pause_setI3028 =>
                \$code_write_request\ <= '0';
                \$v2868\ := eclat_unit;
                \$code_ptr_write\ <= 371;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"11";
                state_var5313 <= pause_setI3027;
              when pause_setI3029 =>
                \$code_write_request\ <= '0';
                \$v2867\ := eclat_unit;
                \$code_ptr_write\ <= 370;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3028;
              when pause_setI3030 =>
                \$code_write_request\ <= '0';
                \$v2866\ := eclat_unit;
                \$code_ptr_write\ <= 369;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"46");
                state_var5313 <= pause_setI3029;
              when pause_setI3031 =>
                \$code_write_request\ <= '0';
                \$v2865\ := eclat_unit;
                \$code_ptr_write\ <= 368;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3030;
              when pause_setI3032 =>
                \$code_write_request\ <= '0';
                \$v2864\ := eclat_unit;
                \$code_ptr_write\ <= 367;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3031;
              when pause_setI3033 =>
                \$code_write_request\ <= '0';
                \$v2863\ := eclat_unit;
                \$code_ptr_write\ <= 366;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"15";
                state_var5313 <= pause_setI3032;
              when pause_setI3034 =>
                \$code_write_request\ <= '0';
                \$v2862\ := eclat_unit;
                \$code_ptr_write\ <= 365;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3033;
              when pause_setI3035 =>
                \$code_write_request\ <= '0';
                \$v2861\ := eclat_unit;
                \$code_ptr_write\ <= 364;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3034;
              when pause_setI3036 =>
                \$code_write_request\ <= '0';
                \$v2860\ := eclat_unit;
                \$code_ptr_write\ <= 363;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"0000" & X"12a");
                state_var5313 <= pause_setI3035;
              when pause_setI3037 =>
                \$code_write_request\ <= '0';
                \$v2859\ := eclat_unit;
                \$code_ptr_write\ <= 362;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3036;
              when pause_setI3038 =>
                \$code_write_request\ <= '0';
                \$v2858\ := eclat_unit;
                \$code_ptr_write\ <= 361;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3037;
              when pause_setI3039 =>
                \$code_write_request\ <= '0';
                \$v2857\ := eclat_unit;
                \$code_ptr_write\ <= 360;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3038;
              when pause_setI3040 =>
                \$code_write_request\ <= '0';
                \$v2856\ := eclat_unit;
                \$code_ptr_write\ <= 359;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"12";
                state_var5313 <= pause_setI3039;
              when pause_setI3041 =>
                \$code_write_request\ <= '0';
                \$v2855\ := eclat_unit;
                \$code_ptr_write\ <= 358;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3040;
              when pause_setI3042 =>
                \$code_write_request\ <= '0';
                \$v2854\ := eclat_unit;
                \$code_ptr_write\ <= 357;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3041;
              when pause_setI3043 =>
                \$code_write_request\ <= '0';
                \$v2853\ := eclat_unit;
                \$code_ptr_write\ <= 356;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"0000" & X"138");
                state_var5313 <= pause_setI3042;
              when pause_setI3044 =>
                \$code_write_request\ <= '0';
                \$v2852\ := eclat_unit;
                \$code_ptr_write\ <= 355;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3043;
              when pause_setI3045 =>
                \$code_write_request\ <= '0';
                \$v2851\ := eclat_unit;
                \$code_ptr_write\ <= 354;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3044;
              when pause_setI3046 =>
                \$code_write_request\ <= '0';
                \$v2850\ := eclat_unit;
                \$code_ptr_write\ <= 353;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3045;
              when pause_setI3047 =>
                \$code_write_request\ <= '0';
                \$v2849\ := eclat_unit;
                \$code_ptr_write\ <= 352;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3046;
              when pause_setI3048 =>
                \$code_write_request\ <= '0';
                \$v2848\ := eclat_unit;
                \$code_ptr_write\ <= 351;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3047;
              when pause_setI3049 =>
                \$code_write_request\ <= '0';
                \$v2847\ := eclat_unit;
                \$code_ptr_write\ <= 350;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"23");
                state_var5313 <= pause_setI3048;
              when pause_setI3050 =>
                \$code_write_request\ <= '0';
                \$v2846\ := eclat_unit;
                \$code_ptr_write\ <= 349;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3049;
              when pause_setI3051 =>
                \$code_write_request\ <= '0';
                \$v2845\ := eclat_unit;
                \$code_ptr_write\ <= 348;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3050;
              when pause_setI3052 =>
                \$code_write_request\ <= '0';
                \$v2844\ := eclat_unit;
                \$code_ptr_write\ <= 347;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"14";
                state_var5313 <= pause_setI3051;
              when pause_setI3053 =>
                \$code_write_request\ <= '0';
                \$v2843\ := eclat_unit;
                \$code_ptr_write\ <= 346;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3052;
              when pause_setI3054 =>
                \$code_write_request\ <= '0';
                \$v2842\ := eclat_unit;
                \$code_ptr_write\ <= 345;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"13");
                state_var5313 <= pause_setI3053;
              when pause_setI3055 =>
                \$code_write_request\ <= '0';
                \$v2841\ := eclat_unit;
                \$code_ptr_write\ <= 344;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3054;
              when pause_setI3056 =>
                \$code_write_request\ <= '0';
                \$v2840\ := eclat_unit;
                \$code_ptr_write\ <= 343;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3055;
              when pause_setI3057 =>
                \$code_write_request\ <= '0';
                \$v2839\ := eclat_unit;
                \$code_ptr_write\ <= 342;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"16";
                state_var5313 <= pause_setI3056;
              when pause_setI3058 =>
                \$code_write_request\ <= '0';
                \$v2838\ := eclat_unit;
                \$code_ptr_write\ <= 341;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"39";
                state_var5313 <= pause_setI3057;
              when pause_setI3059 =>
                \$code_write_request\ <= '0';
                \$v2837\ := eclat_unit;
                \$code_ptr_write\ <= 340;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3058;
              when pause_setI3060 =>
                \$code_write_request\ <= '0';
                \$v2836\ := eclat_unit;
                \$code_ptr_write\ <= 339;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"0000" & X"13a");
                state_var5313 <= pause_setI3059;
              when pause_setI3061 =>
                \$code_write_request\ <= '0';
                \$v2835\ := eclat_unit;
                \$code_ptr_write\ <= 338;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3060;
              when pause_setI3062 =>
                \$code_write_request\ <= '0';
                \$v2834\ := eclat_unit;
                \$code_ptr_write\ <= 337;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3061;
              when pause_setI3063 =>
                \$code_write_request\ <= '0';
                \$v2833\ := eclat_unit;
                \$code_ptr_write\ <= 336;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3062;
              when pause_setI3064 =>
                \$code_write_request\ <= '0';
                \$v2832\ := eclat_unit;
                \$code_ptr_write\ <= 335;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"0000" & X"14c");
                state_var5313 <= pause_setI3063;
              when pause_setI3065 =>
                \$code_write_request\ <= '0';
                \$v2831\ := eclat_unit;
                \$code_ptr_write\ <= 334;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3064;
              when pause_setI3066 =>
                \$code_write_request\ <= '0';
                \$v2830\ := eclat_unit;
                \$code_ptr_write\ <= 333;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3065;
              when pause_setI3067 =>
                \$code_write_request\ <= '0';
                \$v2829\ := eclat_unit;
                \$code_ptr_write\ <= 332;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3066;
              when pause_setI3068 =>
                \$code_write_request\ <= '0';
                \$v2828\ := eclat_unit;
                \$code_ptr_write\ <= 331;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3067;
              when pause_setI3069 =>
                \$code_write_request\ <= '0';
                \$v2827\ := eclat_unit;
                \$code_ptr_write\ <= 330;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"26";
                state_var5313 <= pause_setI3068;
              when pause_setI3070 =>
                \$code_write_request\ <= '0';
                \$v2826\ := eclat_unit;
                \$code_ptr_write\ <= 329;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"16";
                state_var5313 <= pause_setI3069;
              when pause_setI3071 =>
                \$code_write_request\ <= '0';
                \$v2825\ := eclat_unit;
                \$code_ptr_write\ <= 328;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3070;
              when pause_setI3072 =>
                \$code_write_request\ <= '0';
                \$v2824\ := eclat_unit;
                \$code_ptr_write\ <= 327;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3071;
              when pause_setI3073 =>
                \$code_write_request\ <= '0';
                \$v2823\ := eclat_unit;
                \$code_ptr_write\ <= 326;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"63";
                state_var5313 <= pause_setI3072;
              when pause_setI3074 =>
                \$code_write_request\ <= '0';
                \$v2822\ := eclat_unit;
                \$code_ptr_write\ <= 325;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3073;
              when pause_setI3075 =>
                \$code_write_request\ <= '0';
                \$v2821\ := eclat_unit;
                \$code_ptr_write\ <= 324;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3074;
              when pause_setI3076 =>
                \$code_write_request\ <= '0';
                \$v2820\ := eclat_unit;
                \$code_ptr_write\ <= 323;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"14";
                state_var5313 <= pause_setI3075;
              when pause_setI3077 =>
                \$code_write_request\ <= '0';
                \$v2819\ := eclat_unit;
                \$code_ptr_write\ <= 322;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3076;
              when pause_setI3078 =>
                \$code_write_request\ <= '0';
                \$v2818\ := eclat_unit;
                \$code_ptr_write\ <= 321;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"22";
                state_var5313 <= pause_setI3077;
              when pause_setI3079 =>
                \$code_write_request\ <= '0';
                \$v2817\ := eclat_unit;
                \$code_ptr_write\ <= 320;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"16";
                state_var5313 <= pause_setI3078;
              when pause_setI3080 =>
                \$code_write_request\ <= '0';
                \$v2816\ := eclat_unit;
                \$code_ptr_write\ <= 319;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3079;
              when pause_setI3081 =>
                \$code_write_request\ <= '0';
                \$v2815\ := eclat_unit;
                \$code_ptr_write\ <= 318;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3080;
              when pause_setI3082 =>
                \$code_write_request\ <= '0';
                \$v2814\ := eclat_unit;
                \$code_ptr_write\ <= 317;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3081;
              when pause_setI3083 =>
                \$code_write_request\ <= '0';
                \$v2813\ := eclat_unit;
                \$code_ptr_write\ <= 316;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3082;
              when pause_setI3084 =>
                \$code_write_request\ <= '0';
                \$v2812\ := eclat_unit;
                \$code_ptr_write\ <= 315;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3083;
              when pause_setI3085 =>
                \$code_write_request\ <= '0';
                \$v2811\ := eclat_unit;
                \$code_ptr_write\ <= 314;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3084;
              when pause_setI3086 =>
                \$code_write_request\ <= '0';
                \$v2810\ := eclat_unit;
                \$code_ptr_write\ <= 313;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3085;
              when pause_setI3087 =>
                \$code_write_request\ <= '0';
                \$v2809\ := eclat_unit;
                \$code_ptr_write\ <= 312;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3086;
              when pause_setI3088 =>
                \$code_write_request\ <= '0';
                \$v2808\ := eclat_unit;
                \$code_ptr_write\ <= 311;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"64";
                state_var5313 <= pause_setI3087;
              when pause_setI3089 =>
                \$code_write_request\ <= '0';
                \$v2807\ := eclat_unit;
                \$code_ptr_write\ <= 310;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3088;
              when pause_setI3090 =>
                \$code_write_request\ <= '0';
                \$v2806\ := eclat_unit;
                \$code_ptr_write\ <= 309;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"27";
                state_var5313 <= pause_setI3089;
              when pause_setI3091 =>
                \$code_write_request\ <= '0';
                \$v2805\ := eclat_unit;
                \$code_ptr_write\ <= 308;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"15";
                state_var5313 <= pause_setI3090;
              when pause_setI3092 =>
                \$code_write_request\ <= '0';
                \$v2804\ := eclat_unit;
                \$code_ptr_write\ <= 307;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3091;
              when pause_setI3093 =>
                \$code_write_request\ <= '0';
                \$v2803\ := eclat_unit;
                \$code_ptr_write\ <= 306;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"69";
                state_var5313 <= pause_setI3092;
              when pause_setI3094 =>
                \$code_write_request\ <= '0';
                \$v2802\ := eclat_unit;
                \$code_ptr_write\ <= 305;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3093;
              when pause_setI3095 =>
                \$code_write_request\ <= '0';
                \$v2801\ := eclat_unit;
                \$code_ptr_write\ <= 304;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3094;
              when pause_setI3096 =>
                \$code_write_request\ <= '0';
                \$v2800\ := eclat_unit;
                \$code_ptr_write\ <= 303;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3095;
              when pause_setI3097 =>
                \$code_write_request\ <= '0';
                \$v2799\ := eclat_unit;
                \$code_ptr_write\ <= 302;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3096;
              when pause_setI3098 =>
                \$code_write_request\ <= '0';
                \$v2798\ := eclat_unit;
                \$code_ptr_write\ <= 301;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3097;
              when pause_setI3099 =>
                \$code_write_request\ <= '0';
                \$v2797\ := eclat_unit;
                \$code_ptr_write\ <= 300;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3098;
              when pause_setI3100 =>
                \$code_write_request\ <= '0';
                \$v2796\ := eclat_unit;
                \$code_ptr_write\ <= 299;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3099;
              when pause_setI3101 =>
                \$code_write_request\ <= '0';
                \$v2795\ := eclat_unit;
                \$code_ptr_write\ <= 298;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3100;
              when pause_setI3102 =>
                \$code_write_request\ <= '0';
                \$v2794\ := eclat_unit;
                \$code_ptr_write\ <= 297;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3101;
              when pause_setI3103 =>
                \$code_write_request\ <= '0';
                \$v2793\ := eclat_unit;
                \$code_ptr_write\ <= 296;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3102;
              when pause_setI3104 =>
                \$code_write_request\ <= '0';
                \$v2792\ := eclat_unit;
                \$code_ptr_write\ <= 295;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3103;
              when pause_setI3105 =>
                \$code_write_request\ <= '0';
                \$v2791\ := eclat_unit;
                \$code_ptr_write\ <= 294;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3104;
              when pause_setI3106 =>
                \$code_write_request\ <= '0';
                \$v2790\ := eclat_unit;
                \$code_ptr_write\ <= 293;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3105;
              when pause_setI3107 =>
                \$code_write_request\ <= '0';
                \$v2789\ := eclat_unit;
                \$code_ptr_write\ <= 292;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"63";
                state_var5313 <= pause_setI3106;
              when pause_setI3108 =>
                \$code_write_request\ <= '0';
                \$v2788\ := eclat_unit;
                \$code_ptr_write\ <= 291;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"2e");
                state_var5313 <= pause_setI3107;
              when pause_setI3109 =>
                \$code_write_request\ <= '0';
                \$v2787\ := eclat_unit;
                \$code_ptr_write\ <= 290;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3108;
              when pause_setI3110 =>
                \$code_write_request\ <= '0';
                \$v2786\ := eclat_unit;
                \$code_ptr_write\ <= 289;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3109;
              when pause_setI3111 =>
                \$code_write_request\ <= '0';
                \$v2785\ := eclat_unit;
                \$code_ptr_write\ <= 288;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3110;
              when pause_setI3112 =>
                \$code_write_request\ <= '0';
                \$v2784\ := eclat_unit;
                \$code_ptr_write\ <= 287;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"14";
                state_var5313 <= pause_setI3111;
              when pause_setI3113 =>
                \$code_write_request\ <= '0';
                \$v2783\ := eclat_unit;
                \$code_ptr_write\ <= 286;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3112;
              when pause_setI3114 =>
                \$code_write_request\ <= '0';
                \$v2782\ := eclat_unit;
                \$code_ptr_write\ <= 285;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3113;
              when pause_setI3115 =>
                \$code_write_request\ <= '0';
                \$v2781\ := eclat_unit;
                \$code_ptr_write\ <= 284;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3114;
              when pause_setI3116 =>
                \$code_write_request\ <= '0';
                \$v2780\ := eclat_unit;
                \$code_ptr_write\ <= 283;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3115;
              when pause_setI3117 =>
                \$code_write_request\ <= '0';
                \$v2779\ := eclat_unit;
                \$code_ptr_write\ <= 282;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3116;
              when pause_setI3118 =>
                \$code_write_request\ <= '0';
                \$v2778\ := eclat_unit;
                \$code_ptr_write\ <= 281;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3117;
              when pause_setI3119 =>
                \$code_write_request\ <= '0';
                \$v2777\ := eclat_unit;
                \$code_ptr_write\ <= 280;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3118;
              when pause_setI3120 =>
                \$code_write_request\ <= '0';
                \$v2776\ := eclat_unit;
                \$code_ptr_write\ <= 279;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1b";
                state_var5313 <= pause_setI3119;
              when pause_setI3121 =>
                \$code_write_request\ <= '0';
                \$v2775\ := eclat_unit;
                \$code_ptr_write\ <= 278;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3120;
              when pause_setI3122 =>
                \$code_write_request\ <= '0';
                \$v2774\ := eclat_unit;
                \$code_ptr_write\ <= 277;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"6";
                state_var5313 <= pause_setI3121;
              when pause_setI3123 =>
                \$code_write_request\ <= '0';
                \$v2773\ := eclat_unit;
                \$code_ptr_write\ <= 276;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3122;
              when pause_setI3124 =>
                \$code_write_request\ <= '0';
                \$v2772\ := eclat_unit;
                \$code_ptr_write\ <= 275;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3123;
              when pause_setI3125 =>
                \$code_write_request\ <= '0';
                \$v2771\ := eclat_unit;
                \$code_ptr_write\ <= 274;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3124;
              when pause_setI3126 =>
                \$code_write_request\ <= '0';
                \$v2770\ := eclat_unit;
                \$code_ptr_write\ <= 273;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3125;
              when pause_setI3127 =>
                \$code_write_request\ <= '0';
                \$v2769\ := eclat_unit;
                \$code_ptr_write\ <= 272;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3126;
              when pause_setI3128 =>
                \$code_write_request\ <= '0';
                \$v2768\ := eclat_unit;
                \$code_ptr_write\ <= 271;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3127;
              when pause_setI3129 =>
                \$code_write_request\ <= '0';
                \$v2767\ := eclat_unit;
                \$code_ptr_write\ <= 270;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"6";
                state_var5313 <= pause_setI3128;
              when pause_setI3130 =>
                \$code_write_request\ <= '0';
                \$v2766\ := eclat_unit;
                \$code_ptr_write\ <= 269;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3129;
              when pause_setI3131 =>
                \$code_write_request\ <= '0';
                \$v2765\ := eclat_unit;
                \$code_ptr_write\ <= 268;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3130;
              when pause_setI3132 =>
                \$code_write_request\ <= '0';
                \$v2764\ := eclat_unit;
                \$code_ptr_write\ <= 267;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3131;
              when pause_setI3133 =>
                \$code_write_request\ <= '0';
                \$v2763\ := eclat_unit;
                \$code_ptr_write\ <= 266;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3132;
              when pause_setI3134 =>
                \$code_write_request\ <= '0';
                \$v2762\ := eclat_unit;
                \$code_ptr_write\ <= 265;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3133;
              when pause_setI3135 =>
                \$code_write_request\ <= '0';
                \$v2761\ := eclat_unit;
                \$code_ptr_write\ <= 264;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3134;
              when pause_setI3136 =>
                \$code_write_request\ <= '0';
                \$v2760\ := eclat_unit;
                \$code_ptr_write\ <= 263;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3135;
              when pause_setI3137 =>
                \$code_write_request\ <= '0';
                \$v2759\ := eclat_unit;
                \$code_ptr_write\ <= 262;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3136;
              when pause_setI3138 =>
                \$code_write_request\ <= '0';
                \$v2758\ := eclat_unit;
                \$code_ptr_write\ <= 261;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3137;
              when pause_setI3139 =>
                \$code_write_request\ <= '0';
                \$v2757\ := eclat_unit;
                \$code_ptr_write\ <= 260;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3138;
              when pause_setI3140 =>
                \$code_write_request\ <= '0';
                \$v2756\ := eclat_unit;
                \$code_ptr_write\ <= 259;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3139;
              when pause_setI3141 =>
                \$code_write_request\ <= '0';
                \$v2755\ := eclat_unit;
                \$code_ptr_write\ <= 258;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3140;
              when pause_setI3142 =>
                \$code_write_request\ <= '0';
                \$v2754\ := eclat_unit;
                \$code_ptr_write\ <= 257;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1c";
                state_var5313 <= pause_setI3141;
              when pause_setI3143 =>
                \$code_write_request\ <= '0';
                \$v2753\ := eclat_unit;
                \$code_ptr_write\ <= 256;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3142;
              when pause_setI3144 =>
                \$code_write_request\ <= '0';
                \$v2752\ := eclat_unit;
                \$code_ptr_write\ <= 255;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3143;
              when pause_setI3145 =>
                \$code_write_request\ <= '0';
                \$v2751\ := eclat_unit;
                \$code_ptr_write\ <= 254;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3144;
              when pause_setI3146 =>
                \$code_write_request\ <= '0';
                \$v2750\ := eclat_unit;
                \$code_ptr_write\ <= 253;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3145;
              when pause_setI3147 =>
                \$code_write_request\ <= '0';
                \$v2749\ := eclat_unit;
                \$code_ptr_write\ <= 252;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3146;
              when pause_setI3148 =>
                \$code_write_request\ <= '0';
                \$v2748\ := eclat_unit;
                \$code_ptr_write\ <= 251;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1b";
                state_var5313 <= pause_setI3147;
              when pause_setI3149 =>
                \$code_write_request\ <= '0';
                \$v2747\ := eclat_unit;
                \$code_ptr_write\ <= 250;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3148;
              when pause_setI3150 =>
                \$code_write_request\ <= '0';
                \$v2746\ := eclat_unit;
                \$code_ptr_write\ <= 249;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3149;
              when pause_setI3151 =>
                \$code_write_request\ <= '0';
                \$v2745\ := eclat_unit;
                \$code_ptr_write\ <= 248;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3150;
              when pause_setI3152 =>
                \$code_write_request\ <= '0';
                \$v2744\ := eclat_unit;
                \$code_ptr_write\ <= 247;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3151;
              when pause_setI3153 =>
                \$code_write_request\ <= '0';
                \$v2743\ := eclat_unit;
                \$code_ptr_write\ <= 246;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3152;
              when pause_setI3154 =>
                \$code_write_request\ <= '0';
                \$v2742\ := eclat_unit;
                \$code_ptr_write\ <= 245;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3153;
              when pause_setI3155 =>
                \$code_write_request\ <= '0';
                \$v2741\ := eclat_unit;
                \$code_ptr_write\ <= 244;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3154;
              when pause_setI3156 =>
                \$code_write_request\ <= '0';
                \$v2740\ := eclat_unit;
                \$code_ptr_write\ <= 243;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3155;
              when pause_setI3157 =>
                \$code_write_request\ <= '0';
                \$v2739\ := eclat_unit;
                \$code_ptr_write\ <= 242;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3156;
              when pause_setI3158 =>
                \$code_write_request\ <= '0';
                \$v2738\ := eclat_unit;
                \$code_ptr_write\ <= 241;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3157;
              when pause_setI3159 =>
                \$code_write_request\ <= '0';
                \$v2737\ := eclat_unit;
                \$code_ptr_write\ <= 240;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3158;
              when pause_setI3160 =>
                \$code_write_request\ <= '0';
                \$v2736\ := eclat_unit;
                \$code_ptr_write\ <= 239;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3159;
              when pause_setI3161 =>
                \$code_write_request\ <= '0';
                \$v2735\ := eclat_unit;
                \$code_ptr_write\ <= 238;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"63";
                state_var5313 <= pause_setI3160;
              when pause_setI3162 =>
                \$code_write_request\ <= '0';
                \$v2734\ := eclat_unit;
                \$code_ptr_write\ <= 237;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"23");
                state_var5313 <= pause_setI3161;
              when pause_setI3163 =>
                \$code_write_request\ <= '0';
                \$v2733\ := eclat_unit;
                \$code_ptr_write\ <= 236;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3162;
              when pause_setI3164 =>
                \$code_write_request\ <= '0';
                \$v2732\ := eclat_unit;
                \$code_ptr_write\ <= 235;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3163;
              when pause_setI3165 =>
                \$code_write_request\ <= '0';
                \$v2731\ := eclat_unit;
                \$code_ptr_write\ <= 234;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3164;
              when pause_setI3166 =>
                \$code_write_request\ <= '0';
                \$v2730\ := eclat_unit;
                \$code_ptr_write\ <= 233;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"14";
                state_var5313 <= pause_setI3165;
              when pause_setI3167 =>
                \$code_write_request\ <= '0';
                \$v2729\ := eclat_unit;
                \$code_ptr_write\ <= 232;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3166;
              when pause_setI3168 =>
                \$code_write_request\ <= '0';
                \$v2728\ := eclat_unit;
                \$code_ptr_write\ <= 231;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3167;
              when pause_setI3169 =>
                \$code_write_request\ <= '0';
                \$v2727\ := eclat_unit;
                \$code_ptr_write\ <= 230;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3168;
              when pause_setI3170 =>
                \$code_write_request\ <= '0';
                \$v2726\ := eclat_unit;
                \$code_ptr_write\ <= 229;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3169;
              when pause_setI3171 =>
                \$code_write_request\ <= '0';
                \$v2725\ := eclat_unit;
                \$code_ptr_write\ <= 228;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3170;
              when pause_setI3172 =>
                \$code_write_request\ <= '0';
                \$v2724\ := eclat_unit;
                \$code_ptr_write\ <= 227;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3171;
              when pause_setI3173 =>
                \$code_write_request\ <= '0';
                \$v2723\ := eclat_unit;
                \$code_ptr_write\ <= 226;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3172;
              when pause_setI3174 =>
                \$code_write_request\ <= '0';
                \$v2722\ := eclat_unit;
                \$code_ptr_write\ <= 225;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1b";
                state_var5313 <= pause_setI3173;
              when pause_setI3175 =>
                \$code_write_request\ <= '0';
                \$v2721\ := eclat_unit;
                \$code_ptr_write\ <= 224;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3174;
              when pause_setI3176 =>
                \$code_write_request\ <= '0';
                \$v2720\ := eclat_unit;
                \$code_ptr_write\ <= 223;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"5";
                state_var5313 <= pause_setI3175;
              when pause_setI3177 =>
                \$code_write_request\ <= '0';
                \$v2719\ := eclat_unit;
                \$code_ptr_write\ <= 222;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3176;
              when pause_setI3178 =>
                \$code_write_request\ <= '0';
                \$v2718\ := eclat_unit;
                \$code_ptr_write\ <= 221;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3177;
              when pause_setI3179 =>
                \$code_write_request\ <= '0';
                \$v2717\ := eclat_unit;
                \$code_ptr_write\ <= 220;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3178;
              when pause_setI3180 =>
                \$code_write_request\ <= '0';
                \$v2716\ := eclat_unit;
                \$code_ptr_write\ <= 219;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3179;
              when pause_setI3181 =>
                \$code_write_request\ <= '0';
                \$v2715\ := eclat_unit;
                \$code_ptr_write\ <= 218;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3180;
              when pause_setI3182 =>
                \$code_write_request\ <= '0';
                \$v2714\ := eclat_unit;
                \$code_ptr_write\ <= 217;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3181;
              when pause_setI3183 =>
                \$code_write_request\ <= '0';
                \$v2713\ := eclat_unit;
                \$code_ptr_write\ <= 216;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3182;
              when pause_setI3184 =>
                \$code_write_request\ <= '0';
                \$v2712\ := eclat_unit;
                \$code_ptr_write\ <= 215;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3183;
              when pause_setI3185 =>
                \$code_write_request\ <= '0';
                \$v2711\ := eclat_unit;
                \$code_ptr_write\ <= 214;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3184;
              when pause_setI3186 =>
                \$code_write_request\ <= '0';
                \$v2710\ := eclat_unit;
                \$code_ptr_write\ <= 213;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3185;
              when pause_setI3187 =>
                \$code_write_request\ <= '0';
                \$v2709\ := eclat_unit;
                \$code_ptr_write\ <= 212;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3186;
              when pause_setI3188 =>
                \$code_write_request\ <= '0';
                \$v2708\ := eclat_unit;
                \$code_ptr_write\ <= 211;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1c";
                state_var5313 <= pause_setI3187;
              when pause_setI3189 =>
                \$code_write_request\ <= '0';
                \$v2707\ := eclat_unit;
                \$code_ptr_write\ <= 210;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3188;
              when pause_setI3190 =>
                \$code_write_request\ <= '0';
                \$v2706\ := eclat_unit;
                \$code_ptr_write\ <= 209;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3189;
              when pause_setI3191 =>
                \$code_write_request\ <= '0';
                \$v2705\ := eclat_unit;
                \$code_ptr_write\ <= 208;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"10";
                state_var5313 <= pause_setI3190;
              when pause_setI3192 =>
                \$code_write_request\ <= '0';
                \$v2704\ := eclat_unit;
                \$code_ptr_write\ <= 207;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3191;
              when pause_setI3193 =>
                \$code_write_request\ <= '0';
                \$v2703\ := eclat_unit;
                \$code_ptr_write\ <= 206;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3192;
              when pause_setI3194 =>
                \$code_write_request\ <= '0';
                \$v2702\ := eclat_unit;
                \$code_ptr_write\ <= 205;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3193;
              when pause_setI3195 =>
                \$code_write_request\ <= '0';
                \$v2701\ := eclat_unit;
                \$code_ptr_write\ <= 204;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3194;
              when pause_setI3196 =>
                \$code_write_request\ <= '0';
                \$v2700\ := eclat_unit;
                \$code_ptr_write\ <= 203;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3195;
              when pause_setI3197 =>
                \$code_write_request\ <= '0';
                \$v2699\ := eclat_unit;
                \$code_ptr_write\ <= 202;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3196;
              when pause_setI3198 =>
                \$code_write_request\ <= '0';
                \$v2698\ := eclat_unit;
                \$code_ptr_write\ <= 201;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3197;
              when pause_setI3199 =>
                \$code_write_request\ <= '0';
                \$v2697\ := eclat_unit;
                \$code_ptr_write\ <= 200;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3198;
              when pause_setI3200 =>
                \$code_write_request\ <= '0';
                \$v2696\ := eclat_unit;
                \$code_ptr_write\ <= 199;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3199;
              when pause_setI3201 =>
                \$code_write_request\ <= '0';
                \$v2695\ := eclat_unit;
                \$code_ptr_write\ <= 198;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3200;
              when pause_setI3202 =>
                \$code_write_request\ <= '0';
                \$v2694\ := eclat_unit;
                \$code_ptr_write\ <= 197;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3201;
              when pause_setI3203 =>
                \$code_write_request\ <= '0';
                \$v2693\ := eclat_unit;
                \$code_ptr_write\ <= 196;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3202;
              when pause_setI3204 =>
                \$code_write_request\ <= '0';
                \$v2692\ := eclat_unit;
                \$code_ptr_write\ <= 195;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"63";
                state_var5313 <= pause_setI3203;
              when pause_setI3205 =>
                \$code_write_request\ <= '0';
                \$v2691\ := eclat_unit;
                \$code_ptr_write\ <= 194;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"17");
                state_var5313 <= pause_setI3204;
              when pause_setI3206 =>
                \$code_write_request\ <= '0';
                \$v2690\ := eclat_unit;
                \$code_ptr_write\ <= 193;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3205;
              when pause_setI3207 =>
                \$code_write_request\ <= '0';
                \$v2689\ := eclat_unit;
                \$code_ptr_write\ <= 192;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3206;
              when pause_setI3208 =>
                \$code_write_request\ <= '0';
                \$v2688\ := eclat_unit;
                \$code_ptr_write\ <= 191;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3207;
              when pause_setI3209 =>
                \$code_write_request\ <= '0';
                \$v2687\ := eclat_unit;
                \$code_ptr_write\ <= 190;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3208;
              when pause_setI3210 =>
                \$code_write_request\ <= '0';
                \$v2686\ := eclat_unit;
                \$code_ptr_write\ <= 189;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3209;
              when pause_setI3211 =>
                \$code_write_request\ <= '0';
                \$v2685\ := eclat_unit;
                \$code_ptr_write\ <= 188;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3210;
              when pause_setI3212 =>
                \$code_write_request\ <= '0';
                \$v2684\ := eclat_unit;
                \$code_ptr_write\ <= 187;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3211;
              when pause_setI3213 =>
                \$code_write_request\ <= '0';
                \$v2683\ := eclat_unit;
                \$code_ptr_write\ <= 186;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3212;
              when pause_setI3214 =>
                \$code_write_request\ <= '0';
                \$v2682\ := eclat_unit;
                \$code_ptr_write\ <= 185;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3213;
              when pause_setI3215 =>
                \$code_write_request\ <= '0';
                \$v2681\ := eclat_unit;
                \$code_ptr_write\ <= 184;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3214;
              when pause_setI3216 =>
                \$code_write_request\ <= '0';
                \$v2680\ := eclat_unit;
                \$code_ptr_write\ <= 183;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3215;
              when pause_setI3217 =>
                \$code_write_request\ <= '0';
                \$v2679\ := eclat_unit;
                \$code_ptr_write\ <= 182;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3216;
              when pause_setI3218 =>
                \$code_write_request\ <= '0';
                \$v2678\ := eclat_unit;
                \$code_ptr_write\ <= 181;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3217;
              when pause_setI3219 =>
                \$code_write_request\ <= '0';
                \$v2677\ := eclat_unit;
                \$code_ptr_write\ <= 180;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3218;
              when pause_setI3220 =>
                \$code_write_request\ <= '0';
                \$v2676\ := eclat_unit;
                \$code_ptr_write\ <= 179;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7f";
                state_var5313 <= pause_setI3219;
              when pause_setI3221 =>
                \$code_write_request\ <= '0';
                \$v2675\ := eclat_unit;
                \$code_ptr_write\ <= 178;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3220;
              when pause_setI3222 =>
                \$code_write_request\ <= '0';
                \$v2674\ := eclat_unit;
                \$code_ptr_write\ <= 177;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3221;
              when pause_setI3223 =>
                \$code_write_request\ <= '0';
                \$v2673\ := eclat_unit;
                \$code_ptr_write\ <= 176;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3222;
              when pause_setI3224 =>
                \$code_write_request\ <= '0';
                \$v2672\ := eclat_unit;
                \$code_ptr_write\ <= 175;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3223;
              when pause_setI3225 =>
                \$code_write_request\ <= '0';
                \$v2671\ := eclat_unit;
                \$code_ptr_write\ <= 174;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3224;
              when pause_setI3226 =>
                \$code_write_request\ <= '0';
                \$v2670\ := eclat_unit;
                \$code_ptr_write\ <= 173;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3225;
              when pause_setI3227 =>
                \$code_write_request\ <= '0';
                \$v2669\ := eclat_unit;
                \$code_ptr_write\ <= 172;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3226;
              when pause_setI3228 =>
                \$code_write_request\ <= '0';
                \$v2668\ := eclat_unit;
                \$code_ptr_write\ <= 171;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3227;
              when pause_setI3229 =>
                \$code_write_request\ <= '0';
                \$v2667\ := eclat_unit;
                \$code_ptr_write\ <= 170;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"5";
                state_var5313 <= pause_setI3228;
              when pause_setI3230 =>
                \$code_write_request\ <= '0';
                \$v2666\ := eclat_unit;
                \$code_ptr_write\ <= 169;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"25";
                state_var5313 <= pause_setI3229;
              when pause_setI3231 =>
                \$code_write_request\ <= '0';
                \$v2665\ := eclat_unit;
                \$code_ptr_write\ <= 168;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"13";
                state_var5313 <= pause_setI3230;
              when pause_setI3232 =>
                \$code_write_request\ <= '0';
                \$v2664\ := eclat_unit;
                \$code_ptr_write\ <= 167;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3231;
              when pause_setI3233 =>
                \$code_write_request\ <= '0';
                \$v2663\ := eclat_unit;
                \$code_ptr_write\ <= 166;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3232;
              when pause_setI3234 =>
                \$code_write_request\ <= '0';
                \$v2662\ := eclat_unit;
                \$code_ptr_write\ <= 165;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3233;
              when pause_setI3235 =>
                \$code_write_request\ <= '0';
                \$v2661\ := eclat_unit;
                \$code_ptr_write\ <= 164;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3234;
              when pause_setI3236 =>
                \$code_write_request\ <= '0';
                \$v2660\ := eclat_unit;
                \$code_ptr_write\ <= 163;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"37");
                state_var5313 <= pause_setI3235;
              when pause_setI3237 =>
                \$code_write_request\ <= '0';
                \$v2659\ := eclat_unit;
                \$code_ptr_write\ <= 162;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3236;
              when pause_setI3238 =>
                \$code_write_request\ <= '0';
                \$v2658\ := eclat_unit;
                \$code_ptr_write\ <= 161;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3237;
              when pause_setI3239 =>
                \$code_write_request\ <= '0';
                \$v2657\ := eclat_unit;
                \$code_ptr_write\ <= 160;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2c";
                state_var5313 <= pause_setI3238;
              when pause_setI3240 =>
                \$code_write_request\ <= '0';
                \$v2656\ := eclat_unit;
                \$code_ptr_write\ <= 159;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"12";
                state_var5313 <= pause_setI3239;
              when pause_setI3241 =>
                \$code_write_request\ <= '0';
                \$v2655\ := eclat_unit;
                \$code_ptr_write\ <= 158;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3240;
              when pause_setI3242 =>
                \$code_write_request\ <= '0';
                \$v2654\ := eclat_unit;
                \$code_ptr_write\ <= 157;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3241;
              when pause_setI3243 =>
                \$code_write_request\ <= '0';
                \$v2653\ := eclat_unit;
                \$code_ptr_write\ <= 156;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"00000" & X"19");
                state_var5313 <= pause_setI3242;
              when pause_setI3244 =>
                \$code_write_request\ <= '0';
                \$v2652\ := eclat_unit;
                \$code_ptr_write\ <= 155;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3243;
              when pause_setI3245 =>
                \$code_write_request\ <= '0';
                \$v2651\ := eclat_unit;
                \$code_ptr_write\ <= 154;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3244;
              when pause_setI3246 =>
                \$code_write_request\ <= '0';
                \$v2650\ := eclat_unit;
                \$code_ptr_write\ <= 153;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"11";
                state_var5313 <= pause_setI3245;
              when pause_setI3247 =>
                \$code_write_request\ <= '0';
                \$v2649\ := eclat_unit;
                \$code_ptr_write\ <= 152;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3246;
              when pause_setI3248 =>
                \$code_write_request\ <= '0';
                \$v2648\ := eclat_unit;
                \$code_ptr_write\ <= 151;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"10";
                state_var5313 <= pause_setI3247;
              when pause_setI3249 =>
                \$code_write_request\ <= '0';
                \$v2647\ := eclat_unit;
                \$code_ptr_write\ <= 150;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3248;
              when pause_setI3250 =>
                \$code_write_request\ <= '0';
                \$v2646\ := eclat_unit;
                \$code_ptr_write\ <= 149;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"f";
                state_var5313 <= pause_setI3249;
              when pause_setI3251 =>
                \$code_write_request\ <= '0';
                \$v2645\ := eclat_unit;
                \$code_ptr_write\ <= 148;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3250;
              when pause_setI3252 =>
                \$code_write_request\ <= '0';
                \$v2644\ := eclat_unit;
                \$code_ptr_write\ <= 147;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3251;
              when pause_setI3253 =>
                \$code_write_request\ <= '0';
                \$v2643\ := eclat_unit;
                \$code_ptr_write\ <= 146;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3252;
              when pause_setI3254 =>
                \$code_write_request\ <= '0';
                \$v2642\ := eclat_unit;
                \$code_ptr_write\ <= 145;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"e";
                state_var5313 <= pause_setI3253;
              when pause_setI3255 =>
                \$code_write_request\ <= '0';
                \$v2641\ := eclat_unit;
                \$code_ptr_write\ <= 144;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3254;
              when pause_setI3256 =>
                \$code_write_request\ <= '0';
                \$v2640\ := eclat_unit;
                \$code_ptr_write\ <= 143;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3255;
              when pause_setI3257 =>
                \$code_write_request\ <= '0';
                \$v2639\ := eclat_unit;
                \$code_ptr_write\ <= 142;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3256;
              when pause_setI3258 =>
                \$code_write_request\ <= '0';
                \$v2638\ := eclat_unit;
                \$code_ptr_write\ <= 141;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"26";
                state_var5313 <= pause_setI3257;
              when pause_setI3259 =>
                \$code_write_request\ <= '0';
                \$v2637\ := eclat_unit;
                \$code_ptr_write\ <= 140;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1c";
                state_var5313 <= pause_setI3258;
              when pause_setI3260 =>
                \$code_write_request\ <= '0';
                \$v2636\ := eclat_unit;
                \$code_ptr_write\ <= 139;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1b";
                state_var5313 <= pause_setI3259;
              when pause_setI3261 =>
                \$code_write_request\ <= '0';
                \$v2635\ := eclat_unit;
                \$code_ptr_write\ <= 138;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"22";
                state_var5313 <= pause_setI3260;
              when pause_setI3262 =>
                \$code_write_request\ <= '0';
                \$v2634\ := eclat_unit;
                \$code_ptr_write\ <= 137;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1d";
                state_var5313 <= pause_setI3261;
              when pause_setI3263 =>
                \$code_write_request\ <= '0';
                \$v2633\ := eclat_unit;
                \$code_ptr_write\ <= 136;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"b");
                state_var5313 <= pause_setI3262;
              when pause_setI3264 =>
                \$code_write_request\ <= '0';
                \$v2632\ := eclat_unit;
                \$code_ptr_write\ <= 135;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3263;
              when pause_setI3265 =>
                \$code_write_request\ <= '0';
                \$v2631\ := eclat_unit;
                \$code_ptr_write\ <= 134;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2b";
                state_var5313 <= pause_setI3264;
              when pause_setI3266 =>
                \$code_write_request\ <= '0';
                \$v2630\ := eclat_unit;
                \$code_ptr_write\ <= 133;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3265;
              when pause_setI3267 =>
                \$code_write_request\ <= '0';
                \$v2629\ := eclat_unit;
                \$code_ptr_write\ <= 132;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"5";
                state_var5313 <= pause_setI3266;
              when pause_setI3268 =>
                \$code_write_request\ <= '0';
                \$v2628\ := eclat_unit;
                \$code_ptr_write\ <= 131;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"19";
                state_var5313 <= pause_setI3267;
              when pause_setI3269 =>
                \$code_write_request\ <= '0';
                \$v2627\ := eclat_unit;
                \$code_ptr_write\ <= 130;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3268;
              when pause_setI3270 =>
                \$code_write_request\ <= '0';
                \$v2626\ := eclat_unit;
                \$code_ptr_write\ <= 129;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3269;
              when pause_setI3271 =>
                \$code_write_request\ <= '0';
                \$v2625\ := eclat_unit;
                \$code_ptr_write\ <= 128;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3270;
              when pause_setI3272 =>
                \$code_write_request\ <= '0';
                \$v2624\ := eclat_unit;
                \$code_ptr_write\ <= 127;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3271;
              when pause_setI3273 =>
                \$code_write_request\ <= '0';
                \$v2623\ := eclat_unit;
                \$code_ptr_write\ <= 126;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3272;
              when pause_setI3274 =>
                \$code_write_request\ <= '0';
                \$v2622\ := eclat_unit;
                \$code_ptr_write\ <= 125;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"16";
                state_var5313 <= pause_setI3273;
              when pause_setI3275 =>
                \$code_write_request\ <= '0';
                \$v2621\ := eclat_unit;
                \$code_ptr_write\ <= 124;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3274;
              when pause_setI3276 =>
                \$code_write_request\ <= '0';
                \$v2620\ := eclat_unit;
                \$code_ptr_write\ <= 123;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3275;
              when pause_setI3277 =>
                \$code_write_request\ <= '0';
                \$v2619\ := eclat_unit;
                \$code_ptr_write\ <= 122;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3276;
              when pause_setI3278 =>
                \$code_write_request\ <= '0';
                \$v2618\ := eclat_unit;
                \$code_ptr_write\ <= 121;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"35";
                state_var5313 <= pause_setI3277;
              when pause_setI3279 =>
                \$code_write_request\ <= '0';
                \$v2617\ := eclat_unit;
                \$code_ptr_write\ <= 120;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3278;
              when pause_setI3280 =>
                \$code_write_request\ <= '0';
                \$v2616\ := eclat_unit;
                \$code_ptr_write\ <= 119;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"26";
                state_var5313 <= pause_setI3279;
              when pause_setI3281 =>
                \$code_write_request\ <= '0';
                \$v2615\ := eclat_unit;
                \$code_ptr_write\ <= 118;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1b";
                state_var5313 <= pause_setI3280;
              when pause_setI3282 =>
                \$code_write_request\ <= '0';
                \$v2614\ := eclat_unit;
                \$code_ptr_write\ <= 117;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1c";
                state_var5313 <= pause_setI3281;
              when pause_setI3283 =>
                \$code_write_request\ <= '0';
                \$v2613\ := eclat_unit;
                \$code_ptr_write\ <= 116;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3282;
              when pause_setI3284 =>
                \$code_write_request\ <= '0';
                \$v2612\ := eclat_unit;
                \$code_ptr_write\ <= 115;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3283;
              when pause_setI3285 =>
                \$code_write_request\ <= '0';
                \$v2611\ := eclat_unit;
                \$code_ptr_write\ <= 114;
                \$code_write_request\ <= '1';
                \$code_write\ <= eclat_sub("000"& X"000000" & X"0" & "000"& X"000000" & X"1");
                state_var5313 <= pause_setI3284;
              when pause_setI3286 =>
                \$code_write_request\ <= '0';
                \$v2610\ := eclat_unit;
                \$code_ptr_write\ <= 113;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7f";
                state_var5313 <= pause_setI3285;
              when pause_setI3287 =>
                \$code_write_request\ <= '0';
                \$v2609\ := eclat_unit;
                \$code_ptr_write\ <= 112;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3286;
              when pause_setI3288 =>
                \$code_write_request\ <= '0';
                \$v2608\ := eclat_unit;
                \$code_ptr_write\ <= 111;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3287;
              when pause_setI3289 =>
                \$code_write_request\ <= '0';
                \$v2607\ := eclat_unit;
                \$code_ptr_write\ <= 110;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3288;
              when pause_setI3290 =>
                \$code_write_request\ <= '0';
                \$v2606\ := eclat_unit;
                \$code_ptr_write\ <= 109;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"83";
                state_var5313 <= pause_setI3289;
              when pause_setI3291 =>
                \$code_write_request\ <= '0';
                \$v2605\ := eclat_unit;
                \$code_ptr_write\ <= 108;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3290;
              when pause_setI3292 =>
                \$code_write_request\ <= '0';
                \$v2604\ := eclat_unit;
                \$code_ptr_write\ <= 107;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3291;
              when pause_setI3293 =>
                \$code_write_request\ <= '0';
                \$v2603\ := eclat_unit;
                \$code_ptr_write\ <= 106;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3292;
              when pause_setI3294 =>
                \$code_write_request\ <= '0';
                \$v2602\ := eclat_unit;
                \$code_ptr_write\ <= 105;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"64";
                state_var5313 <= pause_setI3293;
              when pause_setI3295 =>
                \$code_write_request\ <= '0';
                \$v2601\ := eclat_unit;
                \$code_ptr_write\ <= 104;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3294;
              when pause_setI3296 =>
                \$code_write_request\ <= '0';
                \$v2600\ := eclat_unit;
                \$code_ptr_write\ <= 103;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3295;
              when pause_setI3297 =>
                \$code_write_request\ <= '0';
                \$v2599\ := eclat_unit;
                \$code_ptr_write\ <= 102;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"7";
                state_var5313 <= pause_setI3296;
              when pause_setI3298 =>
                \$code_write_request\ <= '0';
                \$v2598\ := eclat_unit;
                \$code_ptr_write\ <= 101;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"27";
                state_var5313 <= pause_setI3297;
              when pause_setI3299 =>
                \$code_write_request\ <= '0';
                \$v2597\ := eclat_unit;
                \$code_ptr_write\ <= 100;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3298;
              when pause_setI3300 =>
                \$code_write_request\ <= '0';
                \$v2596\ := eclat_unit;
                \$code_ptr_write\ <= 99;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3299;
              when pause_setI3301 =>
                \$code_write_request\ <= '0';
                \$v2595\ := eclat_unit;
                \$code_ptr_write\ <= 98;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7f";
                state_var5313 <= pause_setI3300;
              when pause_setI3302 =>
                \$code_write_request\ <= '0';
                \$v2594\ := eclat_unit;
                \$code_ptr_write\ <= 97;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3301;
              when pause_setI3303 =>
                \$code_write_request\ <= '0';
                \$v2593\ := eclat_unit;
                \$code_ptr_write\ <= 96;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3302;
              when pause_setI3304 =>
                \$code_write_request\ <= '0';
                \$v2592\ := eclat_unit;
                \$code_ptr_write\ <= 95;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3303;
              when pause_setI3305 =>
                \$code_write_request\ <= '0';
                \$v2591\ := eclat_unit;
                \$code_ptr_write\ <= 94;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"3";
                state_var5313 <= pause_setI3304;
              when pause_setI3306 =>
                \$code_write_request\ <= '0';
                \$v2590\ := eclat_unit;
                \$code_ptr_write\ <= 93;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3305;
              when pause_setI3307 =>
                \$code_write_request\ <= '0';
                \$v2589\ := eclat_unit;
                \$code_ptr_write\ <= 92;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3306;
              when pause_setI3308 =>
                \$code_write_request\ <= '0';
                \$v2588\ := eclat_unit;
                \$code_ptr_write\ <= 91;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"58";
                state_var5313 <= pause_setI3307;
              when pause_setI3309 =>
                \$code_write_request\ <= '0';
                \$v2587\ := eclat_unit;
                \$code_ptr_write\ <= 90;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"79";
                state_var5313 <= pause_setI3308;
              when pause_setI3310 =>
                \$code_write_request\ <= '0';
                \$v2586\ := eclat_unit;
                \$code_ptr_write\ <= 89;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3309;
              when pause_setI3311 =>
                \$code_write_request\ <= '0';
                \$v2585\ := eclat_unit;
                \$code_ptr_write\ <= 88;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"6f";
                state_var5313 <= pause_setI3310;
              when pause_setI3312 =>
                \$code_write_request\ <= '0';
                \$v2584\ := eclat_unit;
                \$code_ptr_write\ <= 87;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3311;
              when pause_setI3313 =>
                \$code_write_request\ <= '0';
                \$v2583\ := eclat_unit;
                \$code_ptr_write\ <= 86;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3312;
              when pause_setI3314 =>
                \$code_write_request\ <= '0';
                \$v2582\ := eclat_unit;
                \$code_ptr_write\ <= 85;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"12";
                state_var5313 <= pause_setI3313;
              when pause_setI3315 =>
                \$code_write_request\ <= '0';
                \$v2581\ := eclat_unit;
                \$code_ptr_write\ <= 84;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3314;
              when pause_setI3316 =>
                \$code_write_request\ <= '0';
                \$v2580\ := eclat_unit;
                \$code_ptr_write\ <= 83;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"58";
                state_var5313 <= pause_setI3315;
              when pause_setI3317 =>
                \$code_write_request\ <= '0';
                \$v2579\ := eclat_unit;
                \$code_ptr_write\ <= 82;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"79";
                state_var5313 <= pause_setI3316;
              when pause_setI3318 =>
                \$code_write_request\ <= '0';
                \$v2578\ := eclat_unit;
                \$code_ptr_write\ <= 81;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3317;
              when pause_setI3319 =>
                \$code_write_request\ <= '0';
                \$v2577\ := eclat_unit;
                \$code_ptr_write\ <= 80;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"6e";
                state_var5313 <= pause_setI3318;
              when pause_setI3320 =>
                \$code_write_request\ <= '0';
                \$v2576\ := eclat_unit;
                \$code_ptr_write\ <= 79;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3319;
              when pause_setI3321 =>
                \$code_write_request\ <= '0';
                \$v2575\ := eclat_unit;
                \$code_ptr_write\ <= 78;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3320;
              when pause_setI3322 =>
                \$code_write_request\ <= '0';
                \$v2574\ := eclat_unit;
                \$code_ptr_write\ <= 77;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"1a";
                state_var5313 <= pause_setI3321;
              when pause_setI3323 =>
                \$code_write_request\ <= '0';
                \$v2573\ := eclat_unit;
                \$code_ptr_write\ <= 76;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3322;
              when pause_setI3324 =>
                \$code_write_request\ <= '0';
                \$v2572\ := eclat_unit;
                \$code_ptr_write\ <= 75;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"58";
                state_var5313 <= pause_setI3323;
              when pause_setI3325 =>
                \$code_write_request\ <= '0';
                \$v2571\ := eclat_unit;
                \$code_ptr_write\ <= 74;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"79";
                state_var5313 <= pause_setI3324;
              when pause_setI3326 =>
                \$code_write_request\ <= '0';
                \$v2570\ := eclat_unit;
                \$code_ptr_write\ <= 73;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"d";
                state_var5313 <= pause_setI3325;
              when pause_setI3327 =>
                \$code_write_request\ <= '0';
                \$v2569\ := eclat_unit;
                \$code_ptr_write\ <= 72;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"a";
                state_var5313 <= pause_setI3326;
              when pause_setI3328 =>
                \$code_write_request\ <= '0';
                \$v2568\ := eclat_unit;
                \$code_ptr_write\ <= 71;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3327;
              when pause_setI3329 =>
                \$code_write_request\ <= '0';
                \$v2567\ := eclat_unit;
                \$code_ptr_write\ <= 70;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3328;
              when pause_setI3330 =>
                \$code_write_request\ <= '0';
                \$v2566\ := eclat_unit;
                \$code_ptr_write\ <= 69;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"24";
                state_var5313 <= pause_setI3329;
              when pause_setI3331 =>
                \$code_write_request\ <= '0';
                \$v2565\ := eclat_unit;
                \$code_ptr_write\ <= 68;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3330;
              when pause_setI3332 =>
                \$code_write_request\ <= '0';
                \$v2564\ := eclat_unit;
                \$code_ptr_write\ <= 67;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3331;
              when pause_setI3333 =>
                \$code_write_request\ <= '0';
                \$v2563\ := eclat_unit;
                \$code_ptr_write\ <= 66;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3332;
              when pause_setI3334 =>
                \$code_write_request\ <= '0';
                \$v2562\ := eclat_unit;
                \$code_ptr_write\ <= 65;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3333;
              when pause_setI3335 =>
                \$code_write_request\ <= '0';
                \$v2561\ := eclat_unit;
                \$code_ptr_write\ <= 64;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3334;
              when pause_setI3336 =>
                \$code_write_request\ <= '0';
                \$v2560\ := eclat_unit;
                \$code_ptr_write\ <= 63;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3335;
              when pause_setI3337 =>
                \$code_write_request\ <= '0';
                \$v2559\ := eclat_unit;
                \$code_ptr_write\ <= 62;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3336;
              when pause_setI3338 =>
                \$code_write_request\ <= '0';
                \$v2558\ := eclat_unit;
                \$code_ptr_write\ <= 61;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3337;
              when pause_setI3339 =>
                \$code_write_request\ <= '0';
                \$v2557\ := eclat_unit;
                \$code_ptr_write\ <= 60;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"26";
                state_var5313 <= pause_setI3338;
              when pause_setI3340 =>
                \$code_write_request\ <= '0';
                \$v2556\ := eclat_unit;
                \$code_ptr_write\ <= 59;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3339;
              when pause_setI3341 =>
                \$code_write_request\ <= '0';
                \$v2555\ := eclat_unit;
                \$code_ptr_write\ <= 58;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"36";
                state_var5313 <= pause_setI3340;
              when pause_setI3342 =>
                \$code_write_request\ <= '0';
                \$v2554\ := eclat_unit;
                \$code_ptr_write\ <= 57;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"21";
                state_var5313 <= pause_setI3341;
              when pause_setI3343 =>
                \$code_write_request\ <= '0';
                \$v2553\ := eclat_unit;
                \$code_ptr_write\ <= 56;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3342;
              when pause_setI3344 =>
                \$code_write_request\ <= '0';
                \$v2552\ := eclat_unit;
                \$code_ptr_write\ <= 55;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3343;
              when pause_setI3345 =>
                \$code_write_request\ <= '0';
                \$v2551\ := eclat_unit;
                \$code_ptr_write\ <= 54;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"c";
                state_var5313 <= pause_setI3344;
              when pause_setI3346 =>
                \$code_write_request\ <= '0';
                \$v2550\ := eclat_unit;
                \$code_ptr_write\ <= 53;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"22";
                state_var5313 <= pause_setI3345;
              when pause_setI3347 =>
                \$code_write_request\ <= '0';
                \$v2549\ := eclat_unit;
                \$code_ptr_write\ <= 52;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3346;
              when pause_setI3348 =>
                \$code_write_request\ <= '0';
                \$v2548\ := eclat_unit;
                \$code_ptr_write\ <= 51;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3347;
              when pause_setI3349 =>
                \$code_write_request\ <= '0';
                \$v2547\ := eclat_unit;
                \$code_ptr_write\ <= 50;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3348;
              when pause_setI3350 =>
                \$code_write_request\ <= '0';
                \$v2546\ := eclat_unit;
                \$code_ptr_write\ <= 49;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3349;
              when pause_setI3351 =>
                \$code_write_request\ <= '0';
                \$v2545\ := eclat_unit;
                \$code_ptr_write\ <= 48;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"e";
                state_var5313 <= pause_setI3350;
              when pause_setI3352 =>
                \$code_write_request\ <= '0';
                \$v2544\ := eclat_unit;
                \$code_ptr_write\ <= 47;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3351;
              when pause_setI3353 =>
                \$code_write_request\ <= '0';
                \$v2543\ := eclat_unit;
                \$code_ptr_write\ <= 46;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3352;
              when pause_setI3354 =>
                \$code_write_request\ <= '0';
                \$v2542\ := eclat_unit;
                \$code_ptr_write\ <= 45;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3353;
              when pause_setI3355 =>
                \$code_write_request\ <= '0';
                \$v2541\ := eclat_unit;
                \$code_ptr_write\ <= 44;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3354;
              when pause_setI3356 =>
                \$code_write_request\ <= '0';
                \$v2540\ := eclat_unit;
                \$code_ptr_write\ <= 43;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3355;
              when pause_setI3357 =>
                \$code_write_request\ <= '0';
                \$v2539\ := eclat_unit;
                \$code_ptr_write\ <= 42;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3356;
              when pause_setI3358 =>
                \$code_write_request\ <= '0';
                \$v2538\ := eclat_unit;
                \$code_ptr_write\ <= 41;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3357;
              when pause_setI3359 =>
                \$code_write_request\ <= '0';
                \$v2537\ := eclat_unit;
                \$code_ptr_write\ <= 40;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3358;
              when pause_setI3360 =>
                \$code_write_request\ <= '0';
                \$v2536\ := eclat_unit;
                \$code_ptr_write\ <= 39;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3359;
              when pause_setI3361 =>
                \$code_write_request\ <= '0';
                \$v2535\ := eclat_unit;
                \$code_ptr_write\ <= 38;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"26";
                state_var5313 <= pause_setI3360;
              when pause_setI3362 =>
                \$code_write_request\ <= '0';
                \$v2534\ := eclat_unit;
                \$code_ptr_write\ <= 37;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3361;
              when pause_setI3363 =>
                \$code_write_request\ <= '0';
                \$v2533\ := eclat_unit;
                \$code_ptr_write\ <= 36;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"44";
                state_var5313 <= pause_setI3362;
              when pause_setI3364 =>
                \$code_write_request\ <= '0';
                \$v2532\ := eclat_unit;
                \$code_ptr_write\ <= 35;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3363;
              when pause_setI3365 =>
                \$code_write_request\ <= '0';
                \$v2531\ := eclat_unit;
                \$code_ptr_write\ <= 34;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3364;
              when pause_setI3366 =>
                \$code_write_request\ <= '0';
                \$v2530\ := eclat_unit;
                \$code_ptr_write\ <= 33;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3365;
              when pause_setI3367 =>
                \$code_write_request\ <= '0';
                \$v2529\ := eclat_unit;
                \$code_ptr_write\ <= 32;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"43";
                state_var5313 <= pause_setI3366;
              when pause_setI3368 =>
                \$code_write_request\ <= '0';
                \$v2528\ := eclat_unit;
                \$code_ptr_write\ <= 31;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3367;
              when pause_setI3369 =>
                \$code_write_request\ <= '0';
                \$v2527\ := eclat_unit;
                \$code_ptr_write\ <= 30;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3368;
              when pause_setI3370 =>
                \$code_write_request\ <= '0';
                \$v2526\ := eclat_unit;
                \$code_ptr_write\ <= 29;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3369;
              when pause_setI3371 =>
                \$code_write_request\ <= '0';
                \$v2525\ := eclat_unit;
                \$code_ptr_write\ <= 28;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3370;
              when pause_setI3372 =>
                \$code_write_request\ <= '0';
                \$v2524\ := eclat_unit;
                \$code_ptr_write\ <= 27;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3371;
              when pause_setI3373 =>
                \$code_write_request\ <= '0';
                \$v2523\ := eclat_unit;
                \$code_ptr_write\ <= 26;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3372;
              when pause_setI3374 =>
                \$code_write_request\ <= '0';
                \$v2522\ := eclat_unit;
                \$code_ptr_write\ <= 25;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3373;
              when pause_setI3375 =>
                \$code_write_request\ <= '0';
                \$v2521\ := eclat_unit;
                \$code_ptr_write\ <= 24;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3374;
              when pause_setI3376 =>
                \$code_write_request\ <= '0';
                \$v2520\ := eclat_unit;
                \$code_ptr_write\ <= 23;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3375;
              when pause_setI3377 =>
                \$code_write_request\ <= '0';
                \$v2519\ := eclat_unit;
                \$code_ptr_write\ <= 22;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3376;
              when pause_setI3378 =>
                \$code_write_request\ <= '0';
                \$v2518\ := eclat_unit;
                \$code_ptr_write\ <= 21;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"0";
                state_var5313 <= pause_setI3377;
              when pause_setI3379 =>
                \$code_write_request\ <= '0';
                \$v2517\ := eclat_unit;
                \$code_ptr_write\ <= 20;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"40";
                state_var5313 <= pause_setI3378;
              when pause_setI3380 =>
                \$code_write_request\ <= '0';
                \$v2516\ := eclat_unit;
                \$code_ptr_write\ <= 19;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3379;
              when pause_setI3381 =>
                \$code_write_request\ <= '0';
                \$v2515\ := eclat_unit;
                \$code_ptr_write\ <= 18;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"22";
                state_var5313 <= pause_setI3380;
              when pause_setI3382 =>
                \$code_write_request\ <= '0';
                \$v2514\ := eclat_unit;
                \$code_ptr_write\ <= 17;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"32";
                state_var5313 <= pause_setI3381;
              when pause_setI3383 =>
                \$code_write_request\ <= '0';
                \$v2513\ := eclat_unit;
                \$code_ptr_write\ <= 16;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3382;
              when pause_setI3384 =>
                \$code_write_request\ <= '0';
                \$v2512\ := eclat_unit;
                \$code_ptr_write\ <= 15;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7f";
                state_var5313 <= pause_setI3383;
              when pause_setI3385 =>
                \$code_write_request\ <= '0';
                \$v2511\ := eclat_unit;
                \$code_ptr_write\ <= 14;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3384;
              when pause_setI3386 =>
                \$code_write_request\ <= '0';
                \$v2510\ := eclat_unit;
                \$code_ptr_write\ <= 13;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3385;
              when pause_setI3387 =>
                \$code_write_request\ <= '0';
                \$v2509\ := eclat_unit;
                \$code_ptr_write\ <= 12;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"2";
                state_var5313 <= pause_setI3386;
              when pause_setI3388 =>
                \$code_write_request\ <= '0';
                \$v2508\ := eclat_unit;
                \$code_ptr_write\ <= 11;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"28";
                state_var5313 <= pause_setI3387;
              when pause_setI3389 =>
                \$code_write_request\ <= '0';
                \$v2507\ := eclat_unit;
                \$code_ptr_write\ <= 10;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"63";
                state_var5313 <= pause_setI3388;
              when pause_setI3390 =>
                \$code_write_request\ <= '0';
                \$v2506\ := eclat_unit;
                \$code_ptr_write\ <= 9;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"4";
                state_var5313 <= pause_setI3389;
              when pause_setI3391 =>
                \$code_write_request\ <= '0';
                \$v2505\ := eclat_unit;
                \$code_ptr_write\ <= 8;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"56";
                state_var5313 <= pause_setI3390;
              when pause_setI3392 =>
                \$code_write_request\ <= '0';
                \$v2504\ := eclat_unit;
                \$code_ptr_write\ <= 7;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"7d";
                state_var5313 <= pause_setI3391;
              when pause_setI3393 =>
                \$code_write_request\ <= '0';
                \$v2503\ := eclat_unit;
                \$code_ptr_write\ <= 6;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"b";
                state_var5313 <= pause_setI3392;
              when pause_setI3394 =>
                \$code_write_request\ <= '0';
                \$v2502\ := eclat_unit;
                \$code_ptr_write\ <= 5;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3393;
              when pause_setI3395 =>
                \$code_write_request\ <= '0';
                \$v2501\ := eclat_unit;
                \$code_ptr_write\ <= 4;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"000000" & X"1";
                state_var5313 <= pause_setI3394;
              when pause_setI3396 =>
                \$code_write_request\ <= '0';
                \$v2500\ := eclat_unit;
                \$code_ptr_write\ <= 3;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"2a";
                state_var5313 <= pause_setI3395;
              when pause_setI3397 =>
                \$code_write_request\ <= '0';
                \$v2499\ := eclat_unit;
                \$code_ptr_write\ <= 2;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"29";
                state_var5313 <= pause_setI3396;
              when pause_setI3398 =>
                \$code_write_request\ <= '0';
                \$v2498\ := eclat_unit;
                \$code_ptr_write\ <= 1;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"0000" & X"14b";
                state_var5313 <= pause_setI3397;
              when pause_setI3399 =>
                \$global_end_write_request\ <= '0';
                \$v2497\ := eclat_unit;
                \$code_ptr_write\ <= 0;
                \$code_write_request\ <= '1';
                \$code_write\ <= "000"& X"00000" & X"54";
                state_var5313 <= pause_setI3398;
              when pause_setI3400 =>
                \$ram_write_request\ <= '0';
                \$v2933\ := eclat_unit;
                \$global_end_ptr_write\ <= 0;
                \$global_end_write_request\ <= '1';
                \$global_end_write\ <= eclat_add(X"3e80" & X"00" & X"17");
                state_var5313 <= pause_setI3399;
              when pause_setI3401 =>
                \$ram_write_request\ <= '0';
                \$v2932\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"16")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3400;
              when pause_setI3402 =>
                \$ram_write_request\ <= '0';
                \$v2931\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"15")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3401;
              when pause_setI3403 =>
                \$ram_write_request\ <= '0';
                \$v2930\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"14")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3402;
              when pause_setI3404 =>
                \$ram_write_request\ <= '0';
                \$v2929\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"13")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3403;
              when pause_setI3405 =>
                \$ram_write_request\ <= '0';
                \$v2928\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"12")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3404;
              when pause_setI3406 =>
                \$ram_write_request\ <= '0';
                \$v2927\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"11")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3405;
              when pause_setI3407 =>
                \$ram_write_request\ <= '0';
                \$v2926\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"00" & X"10")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3406;
              when pause_setI3408 =>
                \$ram_write_request\ <= '0';
                \$v2925\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"f")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3407;
              when pause_setI3409 =>
                \$ram_write_request\ <= '0';
                \$v2924\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"e")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3408;
              when pause_setI3410 =>
                \$ram_write_request\ <= '0';
                \$v2923\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"d")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= eclat_resize(X"3e80",31) & eclat_false;
                state_var5313 <= pause_setI3409;
              when pause_setI3411 =>
                \$ram_write_request\ <= '0';
                \$v2922\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"2")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3410;
              when pause_setI3412 =>
                \$ram_write_request\ <= '0';
                \$v2921\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"1")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3411;
              when pause_setI3413 =>
                \$ram_write_request\ <= '0';
                \$v2920\ := eclat_unit;
                \$ram_ptr_write\ <= 16000;
                \$ram_write_request\ <= '1';
                \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(X"0" & X"0",31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(X"000" & X"2",31) & "000"& X"000000" & X"2")) & eclat_true;
                state_var5313 <= pause_setI3412;
              when compute2976 =>
                rdy2975 := eclat_false;
                \$v1557\ := eclat_unit & eclat_false;
                \$v2496\ := eclat_unit;
                \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & X"000" & X"c")));
                \$ram_write_request\ <= '1';
                \$ram_write\ <= "000"& X"000000" & X"0" & eclat_true;
                state_var5313 <= pause_setI3413;
              end case;
              \$v1824\ := result2974;
              \$v1822\ := \$v1557\;
              \$v1860\ := eclat_not(\$v1556_init\);
              if \$v1860\(0) = '1' then
                \$v1556\ := eclat_false;
                \$v1556_init\ := eclat_true;
              end if;
              \$v1556\ := eclat_and(eclat_if(\$v1556\ & eclat_true & ""&\$v1822\(1)) & eclat_not(eclat_false));
              \$v1823\ := eclat_unit;
              \$548_rdy\ := \$v1556\;
              \$v495\ := eclat_false & eclat_true & \$548_rdy\ & \$v1527\(3 to 10);
              \$v1527\ := \$v495\;
              \$v1810\ := eclat_unit;
              \$v1809\ := \$v1527\;
              \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
              result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
              rdy1858 := eclat_true;
              case compute1859_id is
              when others =>
                
              end case;
            else
              \$v5308\ := eclat_not(\$v1545_init\);
              if \$v5308\(0) = '1' then
                \$v1545\ := X"000" & X"0" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"3e8" & "000"& X"000000" & X"1" & eclat_true & X"0" & X"0" & X"000" & X"0" & eclat_false & eclat_false & eclat_true;
                \$v1545_init\ := eclat_true;
              end if;
              \$v5307\ := eclat_not(""&\$v1527\(2));
              if \$v5307\(0) = '1' then
                \$v232\ := \$v1545\(0 to 121) & eclat_true;
                \$v1545\ := \$v232\;
                \$v1818\ := eclat_unit;
                \$v1814\ := \$v1545\;
                \$v3417\ := ""&\$v1814\(120);
                if \$v3417\(0) = '1' then
                  \$v3416\ := eclat_true;
                  if \$v3416\(0) = '1' then
                    eclat_print_string(of_string("cycle:"));
                    
                    eclat_print_int(\$556_cy\);
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$547_o\ := eclat_false & eclat_true & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false;
                    \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                    \$v1527\ := \$v495\;
                    \$v1810\ := eclat_unit;
                    \$v1809\ := \$v1527\;
                    \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                    result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                    rdy1858 := eclat_true;
                    case compute1859_id is
                    when others =>
                      
                    end case;
                  else
                    \$v1815\ := eclat_unit;
                    \$547_o\ := eclat_false & eclat_true & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false;
                    \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                    \$v1527\ := \$v495\;
                    \$v1810\ := eclat_unit;
                    \$v1809\ := \$v1527\;
                    \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                    result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                    rdy1858 := eclat_true;
                    case compute1859_id is
                    when others =>
                      
                    end case;
                  end if;
                else
                  \$547_o\ := eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_false;
                  \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                  \$v1527\ := \$v495\;
                  \$v1810\ := eclat_unit;
                  \$v1809\ := \$v1527\;
                  \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                  result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                  rdy1858 := eclat_true;
                  case compute1859_id is
                  when others =>
                    
                  end case;
                end if;
              else
                \$v5306\ := eclat_not(\$v1549_init\);
                if \$v5306\(0) = '1' then
                  \$v1549\ := \$v1545\(0 to 121) & eclat_false;
                  \$v1549_init\ := eclat_true;
                end if;
                case state_var5312 is
                when \$706_loop\ =>
                  \$v4924\ := eclat_ge(\$706_loop_arg\(0 to 15) & \$706_loop_arg\(32 to 47));
                  if \$v4924\(0) = '1' then
                    \$706_loop_result\ := eclat_unit;
                    case \$706_loop_id\ is
                    when X"00" & X"1" =>
                      \$v3442\ := \$706_loop_result\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$1603\(0 to 30),16)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$707_copy_root_in_ram_arg\(32 to 47),31) & eclat_false;
                      state_var5312 <= pause_setI4927;
                    when X"00" & X"2" =>
                      \$v3458\ := \$706_loop_result\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$1592\(0 to 30),16)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$708_loop_arg\(16 to 31),31) & eclat_false;
                      state_var5312 <= pause_setI4940;
                    when X"00" & X"7" =>
                      \$v3504\ := \$706_loop_result\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$710_arg\(48 to 78),16)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v3486\(32 to 47),31) & eclat_false;
                      state_var5312 <= pause_setI4958;
                    when X"00" & X"8" =>
                      \$v3517\ := \$706_loop_result\;
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_resize(\$710_arg\(16 to 46),16)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$v3419\(112 to 127),31) & eclat_false;
                      state_var5312 <= pause_setI4967;
                    when others =>
                      
                    end case;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$706_loop_arg\(16 to 31) & \$706_loop_arg\(0 to 15))));
                    state_var5312 <= pause_getI4922;
                  end if;
                when \$707_copy_root_in_ram\ =>
                  \$v4937\ := eclat_ge(\$707_copy_root_in_ram_arg\(0 to 15) & \$707_copy_root_in_ram_arg\(16 to 31));
                  if \$v4937\(0) = '1' then
                    \$707_copy_root_in_ram_result\ := \$707_copy_root_in_ram_arg\(32 to 47);
                    case \$707_copy_root_in_ram_id\ is
                    when X"00" & X"5" =>
                      \$1567_next\ := \$707_copy_root_in_ram_result\;
                      eclat_print_string(of_string("======================================="));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$709_aux_id\ := X"00" & X"4";
                      \$709_aux_arg\ := \$v3419\(112 to 127) & \$1567_next\ & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                      state_var5312 <= \$709_aux\;
                    when X"00" & X"6" =>
                      \$1565_next\ := \$707_copy_root_in_ram_result\;
                      \$global_end_ptr\ <= 0;
                      state_var5312 <= pause_getI4955;
                    when others =>
                      
                    end case;
                  else
                    eclat_print_string(of_string("racine:"));
                    
                    eclat_print_int(\$707_copy_root_in_ram_arg\(0 to 15));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$ram_ptr\ <= to_integer(unsigned(\$707_copy_root_in_ram_arg\(0 to 15)));
                    state_var5312 <= pause_getI4935;
                  end if;
                when \$708_loop\ =>
                  \$v4950\ := eclat_ge(\$708_loop_arg\(0 to 15) & \$708_loop_arg\(32 to 47));
                  if \$v4950\(0) = '1' then
                    \$708_loop_result\ := \$708_loop_arg\(16 to 31);
                    \$1581_next\ := \$708_loop_result\;
                    \$709_aux_arg\ := eclat_add(\$709_aux_arg\(0 to 15) & eclat_add(\$1579\ & X"000" & X"1")) & \$1581_next\ & \$709_aux_arg\(32 to 47) & \$709_aux_arg\(48 to 63) & \$709_aux_arg\(64 to 79);
                    state_var5312 <= \$709_aux\;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(\$708_loop_arg\(80 to 95) & \$708_loop_arg\(0 to 15))));
                    state_var5312 <= pause_getI4948;
                  end if;
                when \$709_aux\ =>
                  eclat_print_string(of_string("     scan="));
                  
                  eclat_print_int(\$709_aux_arg\(0 to 15));
                  
                  eclat_print_string(of_string(" | next="));
                  
                  eclat_print_int(\$709_aux_arg\(16 to 31));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v4953\ := eclat_ge(\$709_aux_arg\(0 to 15) & \$709_aux_arg\(16 to 31));
                  if \$v4953\(0) = '1' then
                    \$709_aux_result\ := \$709_aux_arg\(16 to 31);
                    \$1568_next\ := \$709_aux_result\;
                    eclat_print_string(of_string("memory copied in to_space : "));
                    
                    eclat_print_int(eclat_sub(\$1568_next\ & \$v3419\(112 to 127)));
                    
                    eclat_print_string(of_string(" words"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$v3479\ := \$v3486\(0 to 31) & \$v3487\(0 to 31) & \$1568_next\;
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_string(of_string("[================= GC END ======================]"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$1530\ := \$v3479\(0 to 31) & \$v3479\(32 to 63) & \$v3479\(64 to 79) & eclat_add(\$v3479\(64 to 79) & eclat_add(
                    eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)) & X"000" & X"1")) & \$v3419\(112 to 127) & \$v3419\(96 to 111);
                    \$v3419\ := \$1530\;
                    \$v3478\ := eclat_unit;
                    \$v3477\ := \$v3419\;
                    \$v3468\ := \$v3477\(0 to 31) & \$v3477\(32 to 63) & \$v3477\(64 to 79);
                    eclat_print_string(of_string("size:"));
                    
                    eclat_print_int(eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v3468\(64 to 79)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(\$710_arg\(80 to 87),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(
                    eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)),31) & "000"& X"000000" & X"2")) & eclat_true;
                    state_var5312 <= pause_setI4954;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(\$709_aux_arg\(0 to 15)));
                    state_var5312 <= pause_getI4951;
                  end if;
                when \$710\ =>
                  eclat_print_string(of_string("GC-ALLOC:(size="));
                  
                  eclat_print_int(eclat_add(eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)) & X"000" & X"1"));
                  
                  eclat_print_string(of_string(")"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v4976\ := eclat_not(\$v3419_init\);
                  if \$v4976\(0) = '1' then
                    \$v3419\ := \$710_arg\(16 to 47) & \$710_arg\(48 to 79) & \$710_arg\(120 to 135) & \$710_arg\(120 to 135) & \$710_arg\(120 to 135) & eclat_add(\$710_arg\(120 to 135) & \$710_arg\(104 to 119));
                    \$v3419_init\ := eclat_true;
                  end if;
                  \$v4975\ := eclat_gt(eclat_add(\$v3419\(80 to 95) & eclat_add(
                  eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)) & X"000" & X"1")) & eclat_add(\$v3419\(96 to 111) & \$710_arg\(104 to 119)));
                  if \$v4975\(0) = '1' then
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_string(of_string("[================= GC START ======================]"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$v4974\ := eclat_not(eclat_if(eclat_not(""&\$710_arg\(47)) & 
                                          eclat_if(eclat_le(\$v3419\(96 to 111) & eclat_resize(\$710_arg\(16 to 46),16)) & eclat_lt(eclat_resize(\$710_arg\(16 to 46),16) & eclat_add(\$v3419\(96 to 111) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false));
                    if \$v4974\(0) = '1' then
                      \$v3486\ := \$710_arg\(16 to 47) & \$v3419\(112 to 127);
                      \$v4965\ := eclat_not(eclat_if(eclat_not(""&\$710_arg\(79)) & 
                                            eclat_if(eclat_le(\$v3419\(96 to 111) & eclat_resize(\$710_arg\(48 to 78),16)) & eclat_lt(eclat_resize(\$710_arg\(48 to 78),16) & eclat_add(\$v3419\(96 to 111) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false));
                      if \$v4965\(0) = '1' then
                        \$v3487\ := \$710_arg\(48 to 79) & \$v3486\(32 to 47);
                        \$707_copy_root_in_ram_id\ := X"00" & X"6";
                        \$707_copy_root_in_ram_arg\ := \$710_arg\(152 to 167) & \$710_arg\(0 to 15) & \$v3487\(32 to 47) & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                        state_var5312 <= \$707_copy_root_in_ram\;
                      else
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(48 to 78),16) & X"000" & X"1")));
                        state_var5312 <= pause_getI4963;
                      end if;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(16 to 46),16) & X"000" & X"1")));
                      state_var5312 <= pause_getI4972;
                    end if;
                  else
                    \$1530\ := \$710_arg\(16 to 47) & \$710_arg\(48 to 79) & \$v3419\(80 to 95) & eclat_add(\$v3419\(80 to 95) & eclat_add(
                    eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)) & X"000" & X"1")) & \$v3419\(96 to 111) & \$v3419\(112 to 127);
                    \$v3419\ := \$1530\;
                    \$v3478\ := eclat_unit;
                    \$v3477\ := \$v3419\;
                    \$v3468\ := \$v3477\(0 to 31) & \$v3477\(32 to 63) & \$v3477\(64 to 79);
                    eclat_print_string(of_string("size:"));
                    
                    eclat_print_int(eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v3468\(64 to 79)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_lor(eclat_lsl(eclat_resize(\$710_arg\(80 to 87),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(
                    eclat_if(eclat_eq(\$710_arg\(88 to 103) & X"000" & X"0") & X"000" & X"1" & \$710_arg\(88 to 103)),31) & "000"& X"000000" & X"2")) & eclat_true;
                    state_var5312 <= pause_setI4954;
                  end if;
                when \$711_apply\ =>
                  eclat_print_string(of_string("ENV:"));
                  
                  eclat_print_int(\$711_apply_arg\(92 to 122));
                  
                  eclat_print_string(of_string("<"));
                  
                  \$v4998\ := ""&\$711_apply_arg\(123);
                  if \$v4998\(0) = '1' then
                    eclat_print_string(of_string("int"));
                    
                    eclat_print_string(of_string(">"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$v4997\ := ""&\$711_apply_arg\(0);
                    if \$v4997\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$711_apply_arg\(76 to 91) & X"000" & X"1")));
                      state_var5312 <= pause_getI4995;
                    else
                      \$v3528\ := "000"& X"000000" & X"1" & eclat_true & \$711_apply_arg\(76 to 91);
                      \$v4994\ := ""&\$711_apply_arg\(1);
                      if \$v4994\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3528\(32 to 47) & X"000" & X"1")));
                        state_var5312 <= pause_getI4992;
                      else
                        \$v3529\ := "000"& X"000000" & X"1" & eclat_true & \$v3528\(32 to 47);
                        \$v4991\ := ""&\$711_apply_arg\(2);
                        if \$v4991\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3529\(32 to 47) & X"000" & X"1")));
                          state_var5312 <= pause_getI4989;
                        else
                          \$v3530\ := "000"& X"000000" & X"1" & eclat_true & \$v3529\(32 to 47);
                          \$v4988\ := ""&\$711_apply_arg\(11);
                          if \$v4988\(0) = '1' then
                            \$1275_sp\ := eclat_add(eclat_sub(\$v3530\(32 to 47) & \$711_apply_arg\(12 to 27)) & \$711_apply_arg\(28 to 43));
                            \$v4984\ := ""&\$711_apply_arg\(2);
                            if \$v4984\(0) = '1' then
                              \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$v3530\(0 to 31);
                              state_var5312 <= pause_setI4983;
                            else
                              \$1276_sp\ := \$1275_sp\;
                              \$v4982\ := ""&\$711_apply_arg\(1);
                              if \$v4982\(0) = '1' then
                                \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$v3529\(0 to 31);
                                state_var5312 <= pause_setI4981;
                              else
                                \$1277_sp\ := \$1276_sp\;
                                \$v4980\ := ""&\$711_apply_arg\(0);
                                if \$v4980\(0) = '1' then
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$v3528\(0 to 31);
                                  state_var5312 <= pause_setI4979;
                                else
                                  \$1278_sp\ := \$1277_sp\;
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                                  state_var5312 <= pause_getI4977;
                                end if;
                              end if;
                            end if;
                          else
                            \$ram_ptr_write\ <= to_integer(unsigned(\$v3530\(32 to 47)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(\$711_apply_arg\(124 to 131),31) & eclat_true;
                            state_var5312 <= pause_setI4987;
                          end if;
                        end if;
                      end if;
                    end if;
                  else
                    eclat_print_string(of_string("ptr"));
                    
                    eclat_print_string(of_string(">"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$v4997\ := ""&\$711_apply_arg\(0);
                    if \$v4997\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$711_apply_arg\(76 to 91) & X"000" & X"1")));
                      state_var5312 <= pause_getI4995;
                    else
                      \$v3528\ := "000"& X"000000" & X"1" & eclat_true & \$711_apply_arg\(76 to 91);
                      \$v4994\ := ""&\$711_apply_arg\(1);
                      if \$v4994\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3528\(32 to 47) & X"000" & X"1")));
                        state_var5312 <= pause_getI4992;
                      else
                        \$v3529\ := "000"& X"000000" & X"1" & eclat_true & \$v3528\(32 to 47);
                        \$v4991\ := ""&\$711_apply_arg\(2);
                        if \$v4991\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3529\(32 to 47) & X"000" & X"1")));
                          state_var5312 <= pause_getI4989;
                        else
                          \$v3530\ := "000"& X"000000" & X"1" & eclat_true & \$v3529\(32 to 47);
                          \$v4988\ := ""&\$711_apply_arg\(11);
                          if \$v4988\(0) = '1' then
                            \$1275_sp\ := eclat_add(eclat_sub(\$v3530\(32 to 47) & \$711_apply_arg\(12 to 27)) & \$711_apply_arg\(28 to 43));
                            \$v4984\ := ""&\$711_apply_arg\(2);
                            if \$v4984\(0) = '1' then
                              \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$v3530\(0 to 31);
                              state_var5312 <= pause_setI4983;
                            else
                              \$1276_sp\ := \$1275_sp\;
                              \$v4982\ := ""&\$711_apply_arg\(1);
                              if \$v4982\(0) = '1' then
                                \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                                \$ram_write_request\ <= '1';
                                \$ram_write\ <= \$v3529\(0 to 31);
                                state_var5312 <= pause_setI4981;
                              else
                                \$1277_sp\ := \$1276_sp\;
                                \$v4980\ := ""&\$711_apply_arg\(0);
                                if \$v4980\(0) = '1' then
                                  \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                                  \$ram_write_request\ <= '1';
                                  \$ram_write\ <= \$v3528\(0 to 31);
                                  state_var5312 <= pause_setI4979;
                                else
                                  \$1278_sp\ := \$1277_sp\;
                                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                                  state_var5312 <= pause_getI4977;
                                end if;
                              end if;
                            end if;
                          else
                            \$ram_ptr_write\ <= to_integer(unsigned(\$v3530\(32 to 47)));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= eclat_resize(\$711_apply_arg\(124 to 131),31) & eclat_true;
                            state_var5312 <= pause_setI4987;
                          end if;
                        end if;
                      end if;
                    end if;
                  end if;
                when \$712_offsetclosure_n\ =>
                  \$712_offsetclosure_n_result\ := \$712_offsetclosure_n_arg\(0 to 15) & eclat_resize(eclat_add(eclat_resize(\$712_offsetclosure_n_arg\(48 to 78),16) & \$712_offsetclosure_n_arg\(32 to 47)),31) & eclat_false & \$712_offsetclosure_n_arg\(16 to 31) & \$712_offsetclosure_n_arg\(80 to 135) & \$712_offsetclosure_n_arg\(136 to 137);
                  \$v8\ := \$712_offsetclosure_n_result\;
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when \$713_binop_int\ =>
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$713_binop_int_arg\(65 to 80) & X"000" & X"1")));
                  state_var5312 <= pause_getI5000;
                when \$714_compare\ =>
                  \$v5002\ := \$714_compare_arg\(0 to 31);
                  case \$v5002\ is
                  when X"0000000" & X"0" =>
                    \$714_compare_result\ := eclat_eq(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when X"0000000" & X"1" =>
                    \$714_compare_result\ := eclat_not(eclat_eq(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93)));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when X"0000000" & X"2" =>
                    \$714_compare_result\ := eclat_lt(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when X"0000000" & X"3" =>
                    \$714_compare_result\ := eclat_if(eclat_lt(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93)) & eclat_true & eclat_eq(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93)));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when X"0000000" & X"4" =>
                    \$714_compare_result\ := eclat_not(eclat_if(eclat_lt(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93)) & eclat_true & eclat_eq(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93))));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when X"0000000" & X"5" =>
                    \$714_compare_result\ := eclat_not(eclat_lt(\$714_compare_arg\(32 to 62) & \$714_compare_arg\(63 to 93)));
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  when others =>
                    \$714_compare_result\ := eclat_false;
                    case \$714_compare_id\ is
                    when X"00" & X"9" =>
                      \$1196_res\ := \$714_compare_result\;
                      \$715_binop_compare_result\ := \$715_binop_compare_arg\(138 to 153) & 
                      eclat_if(\$1196_res\ & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v3545\(32 to 47) & \$715_binop_compare_arg\(80 to 135) & \$715_binop_compare_arg\(136 to 137);
                      \$v8\ := \$715_binop_compare_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when X"00" & X"b" =>
                      \$1127_b\ := \$714_compare_result\;
                      \$719_compbranch_result\ := eclat_if(\$1127_b\ & eclat_add(\$719_compbranch_arg\(200 to 215) & eclat_resize(\$719_compbranch_arg\(63 to 93),16)) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199) & \$719_compbranch_arg\(216 to 231) & \$719_compbranch_arg\(94 to 125) & \$719_compbranch_arg\(126 to 141) & \$719_compbranch_arg\(142 to 197) & \$719_compbranch_arg\(198 to 199));
                      \$v8\ := \$719_compbranch_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    when others =>
                      
                    end case;
                  end case;
                when \$715_binop_compare\ =>
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$715_binop_compare_arg\(64 to 79) & X"000" & X"1")));
                  state_var5312 <= pause_getI5003;
                when \$716_make_block_n\ =>
                  \$710_id\ := X"00" & X"a";
                  \$710_arg\ := \$716_make_block_n_arg\(16 to 31) & \$716_make_block_n_arg\(82 to 113) & \$716_make_block_n_arg\(114 to 145) & eclat_resize(\$716_make_block_n_arg\(35 to 65),8) & \$716_make_block_n_arg\(66 to 81) & \$716_make_block_n_arg\(172 to 187) & \$716_make_block_n_arg\(188 to 203) & \$716_make_block_n_arg\(204 to 219) & \$716_make_block_n_arg\(220 to 235);
                  state_var5312 <= \$710\;
                when \$717_branch_if\ =>
                  \$v5017\ := eclat_if(""&\$717_branch_if_arg\(0) & eclat_not(eclat_neq(\$717_branch_if_arg\(1 to 31) & "000"& X"000000" & X"0")) & eclat_neq(\$717_branch_if_arg\(1 to 31) & "000"& X"000000" & X"0"));
                  if \$v5017\(0) = '1' then
                    \$code_ptr\ <= to_integer(unsigned(\$717_branch_if_arg\(107 to 122)));
                    state_var5312 <= pause_getI5015;
                  else
                    \$717_branch_if_result\ := \$717_branch_if_arg\(123 to 138) & \$717_branch_if_arg\(1 to 32) & \$717_branch_if_arg\(33 to 48) & \$717_branch_if_arg\(49 to 104) & \$717_branch_if_arg\(105 to 106);
                    \$v8\ := \$717_branch_if_result\;
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  end if;
                when \$718_loop_push\ =>
                  \$v5021\ := eclat_ge(\$718_loop_push_arg\(16 to 23) & \$718_loop_push_arg\(56 to 63));
                  if \$v5021\(0) = '1' then
                    \$718_loop_push_result\ := \$718_loop_push_arg\(0 to 15);
                    \$970_sp\ := \$718_loop_push_result\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                    state_var5312 <= pause_getI5108;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$718_loop_push_arg\(24 to 54),16) & eclat_resize(eclat_add(\$718_loop_push_arg\(16 to 23) & X"0" & X"2"),16)) & X"000" & X"1")));
                    state_var5312 <= pause_getI5019;
                  end if;
                when \$719_compbranch\ =>
                  \$714_compare_id\ := X"00" & X"b";
                  \$714_compare_arg\ := \$719_compbranch_arg\(0 to 31) & \$719_compbranch_arg\(32 to 62) & \$719_compbranch_arg\(94 to 124);
                  state_var5312 <= \$714_compare\;
                when \$720_w\ =>
                  \$v5025\ := eclat_gt(\$720_w_arg\(0 to 7) & \$720_w_arg\(56 to 63));
                  if \$v5025\(0) = '1' then
                    \$720_w_result\ := \$720_w_arg\(8 to 23);
                    \$859_sp\ := \$720_w_result\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$859_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5199;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$720_w_arg\(8 to 23) & X"000" & X"1")));
                    state_var5312 <= pause_getI5023;
                  end if;
                when \$721_w\ =>
                  \$v5029\ := eclat_gt(\$721_w_arg\(0 to 15) & \$721_w_arg\(32 to 47));
                  if \$v5029\(0) = '1' then
                    \$721_w_result\ := eclat_unit;
                    \$v3594\ := \$721_w_result\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI5270;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$721_w_arg\(16 to 31) & \$721_w_arg\(0 to 15))));
                    state_var5312 <= pause_getI5027;
                  end if;
                when \$722_fill\ =>
                  \$v5033\ := eclat_gt(\$722_fill_arg\(0 to 15) & \$722_fill_arg\(32 to 47));
                  if \$v5033\(0) = '1' then
                    \$722_fill_result\ := \$722_fill_arg\(16 to 31);
                    \$785_sp\ := \$722_fill_result\;
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & \$v3595\(64 to 95) & \$785_sp\ & \$v3595\(32 to 63) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$722_fill_arg\(16 to 31) & X"000" & X"1")));
                    state_var5312 <= pause_getI5031;
                  end if;
                when \$723_fill\ =>
                  \$v5037\ := eclat_ge(\$723_fill_arg\(0 to 15) & \$723_fill_arg\(32 to 47));
                  if \$v5037\(0) = '1' then
                    \$723_fill_result\ := \$723_fill_arg\(16 to 31);
                    \$803_sp\ := \$723_fill_result\;
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & \$v3600\(64 to 95) & \$803_sp\ & \$v3600\(32 to 63) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$723_fill_arg\(16 to 31) & X"000" & X"1")));
                    state_var5312 <= pause_getI5035;
                  end if;
                when \$724_w0\ =>
                  \$v5041\ := eclat_ge(\$724_w0_arg\(0 to 15) & \$724_w0_arg\(32 to 47));
                  if \$v5041\(0) = '1' then
                    \$724_w0_result\ := \$724_w0_arg\(16 to 31);
                    \$762_sp\ := \$724_w0_result\;
                    \$725_w1_id\ := X"0" & X"41";
                    \$725_w1_arg\ := X"000" & X"1" & \$v3589\(64 to 95) & eclat_resize(\$744_argument1\,16) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & X"f9";
                    state_var5312 <= \$725_w1\;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$724_w0_arg\(16 to 31) & X"000" & X"1")));
                    state_var5312 <= pause_getI5039;
                  end if;
                when \$725_w1\ =>
                  \$v5046\ := eclat_ge(\$725_w1_arg\(0 to 15) & \$725_w1_arg\(48 to 63));
                  if \$v5046\(0) = '1' then
                    \$725_w1_result\ := eclat_unit;
                    \$v3591\ := \$725_w1_result\;
                    \$ram_ptr_write\ <= to_integer(unsigned(\$762_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3589\(64 to 95);
                    state_var5312 <= pause_setI5285;
                  else
                    \$1050\ := \$725_w1_arg\(16 to 47) & eclat_sub(eclat_mult(X"000" & X"2" & \$725_w1_arg\(0 to 15)) & X"000" & X"1") & eclat_lor(eclat_lsl(eclat_resize(\$725_w1_arg\(96 to 103),31) & "000"& X"00000" & X"18") & eclat_lsl(eclat_resize(eclat_mult(X"000" & X"2" & \$725_w1_arg\(0 to 15)),31) & "000"& X"000000" & X"2")) & eclat_true;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$1050\(0 to 30),16) & \$1050\(32 to 47)) & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$1050\(48 to 79);
                    state_var5312 <= pause_setI5045;
                  end if;
                when \$726_w3\ =>
                  \$v5048\ := eclat_ge(\$726_w3_arg\(0 to 15) & \$726_w3_arg\(64 to 79));
                  if \$v5048\(0) = '1' then
                    \$726_w3_result\ := \$726_w3_arg\(16 to 31);
                    \$764_sp\ := \$726_w3_result\;
                    \$v8\ := eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & eclat_resize(\$744_argument1\,16)) & \$v3589\(64 to 95) & \$764_sp\ & \$v3589\(32 to 63) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  else
                    \$ram_ptr_write\ <= to_integer(unsigned(\$726_w3_arg\(16 to 31)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(eclat_resize(\$726_w3_arg\(32 to 62),16) & eclat_mult(X"000" & X"2" & \$726_w3_arg\(0 to 15))),31) & eclat_true;
                    state_var5312 <= pause_setI5047;
                  end if;
                when pause_getI5049 =>
                  state_var5312 <= pause_getII5050;
                when pause_getI5051 =>
                  state_var5312 <= pause_getII5052;
                when pause_getI5053 =>
                  state_var5312 <= pause_getII5054;
                when pause_getI5055 =>
                  state_var5312 <= pause_getII5056;
                when pause_getI5057 =>
                  state_var5312 <= pause_getII5058;
                when pause_getI5059 =>
                  state_var5312 <= pause_getII5060;
                when pause_getI5061 =>
                  state_var5312 <= pause_getII5062;
                when pause_getI5063 =>
                  state_var5312 <= pause_getII5064;
                when pause_getI5067 =>
                  state_var5312 <= pause_getII5068;
                when pause_getI5070 =>
                  state_var5312 <= pause_getII5071;
                when pause_getI5073 =>
                  state_var5312 <= pause_getII5074;
                when pause_getI5076 =>
                  state_var5312 <= pause_getII5077;
                when pause_getI5079 =>
                  state_var5312 <= pause_getII5080;
                when pause_getI5082 =>
                  state_var5312 <= pause_getII5083;
                when pause_getI5085 =>
                  state_var5312 <= pause_getII5086;
                when pause_getI5088 =>
                  state_var5312 <= pause_getII5089;
                when pause_getI5090 =>
                  state_var5312 <= pause_getII5091;
                when pause_getI5092 =>
                  state_var5312 <= pause_getII5093;
                when pause_getI5094 =>
                  state_var5312 <= pause_getII5095;
                when pause_getI5096 =>
                  state_var5312 <= pause_getII5097;
                when pause_getI5099 =>
                  state_var5312 <= pause_getII5100;
                when pause_getI5102 =>
                  state_var5312 <= pause_getII5103;
                when pause_getI5105 =>
                  state_var5312 <= pause_getII5106;
                when pause_getI5108 =>
                  state_var5312 <= pause_getII5109;
                when pause_getI5110 =>
                  state_var5312 <= pause_getII5111;
                when pause_getI5116 =>
                  state_var5312 <= pause_getII5117;
                when pause_getI5118 =>
                  state_var5312 <= pause_getII5119;
                when pause_getI5120 =>
                  state_var5312 <= pause_getII5121;
                when pause_getI5122 =>
                  state_var5312 <= pause_getII5123;
                when pause_getI5125 =>
                  state_var5312 <= pause_getII5126;
                when pause_getI5128 =>
                  state_var5312 <= pause_getII5129;
                when pause_getI5131 =>
                  state_var5312 <= pause_getII5132;
                when pause_getI5134 =>
                  state_var5312 <= pause_getII5135;
                when pause_getI5136 =>
                  state_var5312 <= pause_getII5137;
                when pause_getI5138 =>
                  state_var5312 <= pause_getII5139;
                when pause_getI5140 =>
                  state_var5312 <= pause_getII5141;
                when pause_getI5143 =>
                  state_var5312 <= pause_getII5144;
                when pause_getI5145 =>
                  state_var5312 <= pause_getII5146;
                when pause_getI5147 =>
                  state_var5312 <= pause_getII5148;
                when pause_getI5149 =>
                  state_var5312 <= pause_getII5150;
                when pause_getI5152 =>
                  state_var5312 <= pause_getII5153;
                when pause_getI5154 =>
                  state_var5312 <= pause_getII5155;
                when pause_getI5156 =>
                  state_var5312 <= pause_getII5157;
                when pause_getI5158 =>
                  state_var5312 <= pause_getII5159;
                when pause_getI5160 =>
                  state_var5312 <= pause_getII5161;
                when pause_getI5162 =>
                  state_var5312 <= pause_getII5163;
                when pause_getI5164 =>
                  state_var5312 <= pause_getII5165;
                when pause_getI5170 =>
                  state_var5312 <= pause_getII5171;
                when pause_getI5172 =>
                  state_var5312 <= pause_getII5173;
                when pause_getI5176 =>
                  state_var5312 <= pause_getII5177;
                when pause_getI5178 =>
                  state_var5312 <= pause_getII5179;
                when pause_getI5184 =>
                  state_var5312 <= pause_getII5185;
                when pause_getI5186 =>
                  state_var5312 <= pause_getII5187;
                when pause_getI5188 =>
                  state_var5312 <= pause_getII5189;
                when pause_getI5190 =>
                  state_var5312 <= pause_getII5191;
                when pause_getI5192 =>
                  state_var5312 <= pause_getII5193;
                when pause_getI5195 =>
                  state_var5312 <= pause_getII5196;
                when pause_getI5197 =>
                  state_var5312 <= pause_getII5198;
                when pause_getI5199 =>
                  state_var5312 <= pause_getII5200;
                when pause_getI5205 =>
                  state_var5312 <= pause_getII5206;
                when pause_getI5207 =>
                  state_var5312 <= pause_getII5208;
                when pause_getI5212 =>
                  state_var5312 <= pause_getII5213;
                when pause_getI5215 =>
                  state_var5312 <= pause_getII5216;
                when pause_getI5217 =>
                  state_var5312 <= pause_getII5218;
                when pause_getI5219 =>
                  state_var5312 <= pause_getII5220;
                when pause_getI5226 =>
                  state_var5312 <= pause_getII5227;
                when pause_getI5230 =>
                  state_var5312 <= pause_getII5231;
                when pause_getI5234 =>
                  state_var5312 <= pause_getII5235;
                when pause_getI5236 =>
                  state_var5312 <= pause_getII5237;
                when pause_getI5240 =>
                  state_var5312 <= pause_getII5241;
                when pause_getI5242 =>
                  state_var5312 <= pause_getII5243;
                when pause_getI5244 =>
                  state_var5312 <= pause_getII5245;
                when pause_getI5248 =>
                  state_var5312 <= pause_getII5249;
                when pause_getI5250 =>
                  state_var5312 <= pause_getII5251;
                when pause_getI5252 =>
                  state_var5312 <= pause_getII5253;
                when pause_getI5254 =>
                  state_var5312 <= pause_getII5255;
                when pause_getI5258 =>
                  state_var5312 <= pause_getII5259;
                when pause_getI5260 =>
                  state_var5312 <= pause_getII5261;
                when pause_getI5262 =>
                  state_var5312 <= pause_getII5263;
                when pause_getI5264 =>
                  state_var5312 <= pause_getII5265;
                when pause_getI5268 =>
                  state_var5312 <= pause_getII5269;
                when pause_getI5270 =>
                  state_var5312 <= pause_getII5271;
                when pause_getI5275 =>
                  state_var5312 <= pause_getII5276;
                when pause_getI5277 =>
                  state_var5312 <= pause_getII5278;
                when pause_getI5279 =>
                  state_var5312 <= pause_getII5280;
                when pause_getI5281 =>
                  state_var5312 <= pause_getII5282;
                when pause_getI5289 =>
                  state_var5312 <= pause_getII5290;
                when pause_getI5292 =>
                  state_var5312 <= pause_getII5293;
                when pause_getI5295 =>
                  state_var5312 <= pause_getII5296;
                when pause_getI5298 =>
                  state_var5312 <= pause_getII5299;
                when pause_getI5301 =>
                  state_var5312 <= pause_getII5302;
                when pause_getII5050 =>
                  \$5345_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5345_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5052 =>
                  \$5348_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5348_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5054 =>
                  \$5351_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5351_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5056 =>
                  \$5354_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5354_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5058 =>
                  \$5357_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5357_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5060 =>
                  \$5360_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5360_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5062 =>
                  \$5363_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5363_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5064 =>
                  \$5366_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5366_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5068 =>
                  \$5373_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5373_v\ & \$5372_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5071 =>
                  \$5378_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5378_v\ & \$5377_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5074 =>
                  \$5383_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5383_v\ & \$5382_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5077 =>
                  \$5388_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5388_v\ & \$5387_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5080 =>
                  \$5393_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5393_v\ & \$5392_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5083 =>
                  \$5398_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5398_v\ & \$5397_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5086 =>
                  \$5403_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5403_v\ & \$5402_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5089 =>
                  \$5408\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5408\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5091 =>
                  \$5413\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5413\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5093 =>
                  \$5418\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5418\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5095 =>
                  \$5423\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5423\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5097 =>
                  \$5429\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5429\ & \$5427_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5100 =>
                  \$5436\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5436\ & \$5434_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5103 =>
                  \$5443\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5443\ & \$5441_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5106 =>
                  \$5450\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5450\ & \$5448_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5109 =>
                  \$971_next_env\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(16 to 47) & \$970_sp\ & \$971_next_env\ & eclat_add(\$v1545\(96 to 103) & eclat_sub(eclat_resize(\$967\,8) & X"0" & X"2")) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5111 =>
                  \$1667_hd\ := \$ram_value\;
                  \$967\ := eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$1667_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                  \$718_loop_push_id\ := X"00" & X"f";
                  \$718_loop_push_arg\ := \$v1545\(48 to 63) & X"0" & X"0" & \$v1545\(64 to 95) & eclat_sub(eclat_resize(\$967\,8) & X"0" & X"2");
                  state_var5312 <= \$718_loop_push\;
                when pause_getII5117 =>
                  \$5467_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5467_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5119 =>
                  \$5472_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5472_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5121 =>
                  \$5477_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5477_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5123 =>
                  \$5482_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5482_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5126 =>
                  \$5492_v\ := \$ram_value\;
                  \$v3681\ := \$5492_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3681\(0 to 31);
                  state_var5312 <= pause_setI5124;
                when pause_getII5129 =>
                  \$5499_v\ := \$ram_value\;
                  \$v3683\ := \$5499_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3683\(0 to 31);
                  state_var5312 <= pause_setI5127;
                when pause_getII5132 =>
                  \$5506_v\ := \$ram_value\;
                  \$v3685\ := \$5506_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3685\(0 to 31);
                  state_var5312 <= pause_setI5130;
                when pause_getII5135 =>
                  \$5513_v\ := \$ram_value\;
                  \$v3687\ := \$5513_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3687\(0 to 31);
                  state_var5312 <= pause_setI5133;
                when pause_getII5137 =>
                  \$5515_hd\ := \$ram_value\;
                  \$976\ := eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$5515_hd\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_resize(\$976\,31) & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5139 =>
                  \$983_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$983_v\ & \$v3689\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5141 =>
                  \$5523_v\ := \$ram_value\;
                  \$v3689\ := \$5523_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$v3689\(0 to 30),16)) & X"000" & X"1")));
                  state_var5312 <= pause_getI5138;
                when pause_getII5144 =>
                  \$5528_v\ := \$ram_value\;
                  \$v3691\ := \$5528_v\ & eclat_sub(\$v3690\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$v3690\(0 to 30),16)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3691\(0 to 31);
                  state_var5312 <= pause_setI5142;
                when pause_getII5146 =>
                  \$5530_v\ := \$ram_value\;
                  \$v3690\ := \$5530_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3690\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5143;
                when pause_getII5148 =>
                  \$994_next_acc\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$994_next_acc\ & \$v3693\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5150 =>
                  \$5535_v\ := \$ram_value\;
                  \$v3693\ := \$5535_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$v3693\(0 to 30),16)) & X"000" & X"1")));
                  state_var5312 <= pause_getI5147;
                when pause_getII5153 =>
                  \$5540_v\ := \$ram_value\;
                  \$v3695\ := \$5540_v\ & eclat_sub(\$v3694\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$v3694\(0 to 30),16)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3695\(0 to 31);
                  state_var5312 <= pause_setI5151;
                when pause_getII5155 =>
                  \$5542_v\ := \$ram_value\;
                  \$v3694\ := \$5542_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3694\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5152;
                when pause_getII5157 =>
                  \$5544_v\ := \$ram_value\;
                  \$v3697\ := \$5544_v\ & eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1") & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(16 to 47) & eclat_sub(\$v3697\(32 to 47) & X"000" & X"2") & \$v1545\(64 to 95) & \$v1545\(96 to 103) & eclat_resize(\$v3697\(0 to 30),16) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5159 =>
                  \$5546_v\ := \$ram_value\;
                  \$v3701\ := \$5546_v\ & eclat_sub(\$v3700\(32 to 47) & X"000" & X"1");
                  \$v8\ := eclat_resize(\$v3698\(0 to 30),16) & \$v1545\(16 to 47) & \$v3701\(32 to 47) & \$v3700\(0 to 31) & eclat_resize(\$v3701\(0 to 30),8) & eclat_resize(\$v3699\(0 to 30),16) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5161 =>
                  \$5548_v\ := \$ram_value\;
                  \$v3700\ := \$5548_v\ & eclat_sub(\$v3699\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3700\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5158;
                when pause_getII5163 =>
                  \$5550_v\ := \$ram_value\;
                  \$v3699\ := \$5550_v\ & eclat_sub(\$v3698\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3699\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5160;
                when pause_getII5165 =>
                  \$5552_v\ := \$ram_value\;
                  \$v3698\ := \$5552_v\ & eclat_sub(\$v1545\(104 to 119) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3698\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5162;
                when pause_getII5171 =>
                  \$1338_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$1338_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5173 =>
                  \$5243_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$5243_v\ & \$1312_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5177 =>
                  \$1326\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$1326\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5179 =>
                  \$5251\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$5251\ & \$1305_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5185 =>
                  \$821\ := \$ram_value\;
                  \$v8\ := eclat_resize(\$821\(0 to 30),16) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(16 to 47) & eclat_sub(eclat_resize(\$744_argument1\,8) & X"0" & X"1") & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5187 =>
                  \$846\ := \$ram_value\;
                  \$v8\ := eclat_resize(\$846\(0 to 30),16) & \$v1545\(16 to 47) & eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & \$v1545\(16 to 47) & eclat_sub(\$v1545\(96 to 103) & X"0" & X"1") & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5189 =>
                  \$5263_v\ := \$ram_value\;
                  \$v3610\ := \$5263_v\ & eclat_sub(\$v3609\(32 to 47) & X"000" & X"1");
                  \$v8\ := eclat_resize(\$v3608\(0 to 30),16) & \$v1545\(16 to 47) & \$v3610\(32 to 47) & \$v3609\(0 to 31) & eclat_resize(\$v3610\(0 to 30),8) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5191 =>
                  \$5265_v\ := \$ram_value\;
                  \$v3609\ := \$5265_v\ & eclat_sub(\$v3608\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3609\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5188;
                when pause_getII5193 =>
                  \$5267_v\ := \$ram_value\;
                  \$v3608\ := \$5267_v\ & eclat_sub(eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3608\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5190;
                when pause_getII5196 =>
                  \$5272_v\ := \$ram_value\;
                  \$v3616\ := \$5272_v\ & eclat_sub(\$v3615\(32 to 47) & X"000" & X"1");
                  \$v8\ := eclat_resize(\$v3614\(0 to 30),16) & \$v3611\(64 to 95) & \$v3616\(32 to 47) & \$v3615\(0 to 31) & eclat_resize(\$v3616\(0 to 30),8) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5198 =>
                  \$5274_v\ := \$ram_value\;
                  \$v3615\ := \$5274_v\ & eclat_sub(\$v3614\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3615\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5195;
                when pause_getII5200 =>
                  \$5276_v\ := \$ram_value\;
                  \$v3614\ := \$5276_v\ & eclat_sub(\$859_sp\ & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3614\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5197;
                when pause_getII5206 =>
                  \$874_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$874_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5208 =>
                  \$877_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$877_v\ & eclat_add(\$v1545\(48 to 63) & X"000" & X"1") & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5213 =>
                  \$1235_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$1235_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5216 =>
                  \$5295_v\ := \$ram_value\;
                  \$v3622\ := \$5295_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$744_argument1\,16)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3622\(0 to 31);
                  state_var5312 <= pause_setI5214;
                when pause_getII5218 =>
                  \$885\ := \$code_value\;
                  \$v8\ := eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_resize(\$885\,16)) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5220 =>
                  \$1663_hd\ := \$ram_value\;
                  \$888_idx\ := eclat_lsr(eclat_resize(\$1663_hd\(0 to 30),16) & X"00" & X"18");
                  \$883_ofs\ := eclat_add(eclat_resize(\$744_argument1\,16) & \$888_idx\);
                  \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$883_ofs\)));
                  state_var5312 <= pause_getI5217;
                when pause_getII5227 =>
                  \$5303_v\ := \$ram_value\;
                  \$v3629\ := \$5303_v\ & eclat_sub(\$903_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v3628\(0 to 31) & \$v3629\(32 to 47) & \$v3629\(0 to 31) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5231 =>
                  \$5306_v\ := \$ram_value\;
                  \$v3634\ := \$5306_v\ & eclat_sub(\$912_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v3633\(0 to 31) & \$v3634\(32 to 47) & \$v3634\(0 to 31) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5235 =>
                  \$5309_v\ := \$ram_value\;
                  \$v3632\ := \$5309_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3632\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5233;
                when pause_getII5237 =>
                  \$5311_v\ := \$ram_value\;
                  \$v3640\ := \$5311_v\ & eclat_sub(\$923_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v3639\(0 to 31) & \$v3640\(32 to 47) & \$v3640\(0 to 31) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5241 =>
                  \$5314_v\ := \$ram_value\;
                  \$v3638\ := \$5314_v\ & eclat_sub(\$v3637\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3638\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5239;
                when pause_getII5243 =>
                  \$5316_v\ := \$ram_value\;
                  \$v3637\ := \$5316_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3637\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5240;
                when pause_getII5245 =>
                  \$5318_v\ := \$ram_value\;
                  \$v3647\ := \$5318_v\ & eclat_sub(\$936_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v3646\(0 to 31) & \$v3647\(32 to 47) & \$v3647\(0 to 31) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5249 =>
                  \$5321_v\ := \$ram_value\;
                  \$v3645\ := \$5321_v\ & eclat_sub(\$v3644\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3645\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5247;
                when pause_getII5251 =>
                  \$5323_v\ := \$ram_value\;
                  \$v3644\ := \$5323_v\ & eclat_sub(\$v3643\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3644\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5248;
                when pause_getII5253 =>
                  \$5325_v\ := \$ram_value\;
                  \$v3643\ := \$5325_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3643\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5250;
                when pause_getII5255 =>
                  \$5327_v\ := \$ram_value\;
                  \$v3655\ := \$5327_v\ & eclat_sub(\$951_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v3654\(0 to 31) & \$v3655\(32 to 47) & \$v3655\(0 to 31) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5259 =>
                  \$5330_v\ := \$ram_value\;
                  \$v3653\ := \$5330_v\ & eclat_sub(\$v3652\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3653\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5257;
                when pause_getII5261 =>
                  \$5332_v\ := \$ram_value\;
                  \$v3652\ := \$5332_v\ & eclat_sub(\$v3651\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3652\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5258;
                when pause_getII5263 =>
                  \$5334_v\ := \$ram_value\;
                  \$v3651\ := \$5334_v\ & eclat_sub(\$v3650\(32 to 47) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3651\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5260;
                when pause_getII5265 =>
                  \$5336_v\ := \$ram_value\;
                  \$v3650\ := \$5336_v\ & eclat_sub(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3650\(32 to 47) & X"000" & X"1")));
                  state_var5312 <= pause_getI5262;
                when pause_getII5269 =>
                  \$961_f0\ := \$ram_value\;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_add(\$961_f0\(0 to 30) & \$744_argument1\) & eclat_true;
                  state_var5312 <= pause_setI5267;
                when pause_getII5271 =>
                  \$771\ := \$ram_value\;
                  \$v8\ := eclat_resize(\$771\(0 to 30),16) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(16 to 47) & eclat_sub(eclat_add(\$v1545\(96 to 103) & eclat_resize(\$744_argument1\,8)) & X"0" & X"1") & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5276 =>
                  \$790_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & \$790_v\ & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5278 =>
                  \$788\ := \$ram_value\;
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$788\(0 to 30),16) & eclat_resize(\$745_argument2\,16)) & X"000" & X"1")));
                  state_var5312 <= pause_getI5275;
                when pause_getII5280 =>
                  \$796_v\ := \$ram_value\;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & \$796_v\ & eclat_add(\$v1545\(48 to 63) & X"000" & X"1") & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5282 =>
                  \$794\ := \$ram_value\;
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$794\(0 to 30),16) & eclat_resize(\$745_argument2\,16)) & X"000" & X"1")));
                  state_var5312 <= pause_getI5279;
                when pause_getII5290 =>
                  \$747\ := \$code_value\;
                  eclat_print_int(\$747\);
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v8\ := \$v1545\(0 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII5293 =>
                  \$746_argument3\ := \$code_value\;
                  \$v5291\ := eclat_resize(\$740\,8);
                  case \$v5291\ is
                  when X"2c" =>
                    \$v5288\ := eclat_gt(eclat_resize(\$745_argument2\,16) & X"000" & X"0");
                    if \$v5288\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v1545\(16 to 47);
                      state_var5312 <= pause_setI5287;
                    else
                      \$752_sp\ := \$v1545\(48 to 63);
                      \$710_id\ := X"0" & X"43";
                      \$710_arg\ := \$752_sp\ & \$v1545\(16 to 47) & \$v1545\(64 to 95) & X"f7" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(\$744_argument1\,16)) & X"000" & X"1") & eclat_resize(\$745_argument2\,16)) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                      state_var5312 <= \$710\;
                    end if;
                  when others =>
                    eclat_print_string(of_string("unknown opcode : "));
                    
                    \$code_ptr\ <= to_integer(unsigned(\$v1545\(0 to 15)));
                    state_var5312 <= pause_getI5289;
                  end case;
                when pause_getII5296 =>
                  \$745_argument2\ := \$code_value\;
                  \$v5294\ := eclat_resize(\$740\,8);
                  case \$v5294\ is
                  when X"24" =>
                    \$721_w_id\ := X"0" & X"35";
                    \$721_w_arg\ := X"000" & X"1" & \$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16) & eclat_sub(eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & eclat_resize(\$745_argument2\,16));
                    state_var5312 <= \$721_w\;
                  when X"2b" =>
                    \$v5274\ := eclat_gt(eclat_resize(\$744_argument1\,16) & X"000" & X"0");
                    if \$v5274\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v1545\(16 to 47);
                      state_var5312 <= pause_setI5273;
                    else
                      \$778_sp\ := \$v1545\(48 to 63);
                      \$710_id\ := X"0" & X"37";
                      \$710_arg\ := \$778_sp\ & \$v1545\(16 to 47) & \$v1545\(64 to 95) & X"f7" & eclat_add(eclat_resize(\$744_argument1\,16) & X"000" & X"1") & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                      state_var5312 <= \$710\;
                    end if;
                  when X"37" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$744_argument1\,16))));
                    state_var5312 <= pause_getI5277;
                  when X"38" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5283;
                  when X"3e" =>
                    \$710_id\ := X"0" & X"39";
                    \$710_arg\ := \$v1545\(48 to 63) & \$v1545\(16 to 47) & \$v1545\(64 to 95) & eclat_resize(\$745_argument2\,8) & eclat_resize(\$744_argument1\,16) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$710\;
                  when X"83" =>
                    \$719_compbranch_id\ := X"0" & X"3a";
                    \$719_compbranch_arg\ := X"0000000" & X"0" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"84" =>
                    \$719_compbranch_id\ := X"0" & X"3b";
                    \$719_compbranch_arg\ := X"0000000" & X"1" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"85" =>
                    \$719_compbranch_id\ := X"0" & X"3c";
                    \$719_compbranch_arg\ := X"0000000" & X"2" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"86" =>
                    \$719_compbranch_id\ := X"0" & X"3d";
                    \$719_compbranch_arg\ := X"0000000" & X"3" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"87" =>
                    \$719_compbranch_id\ := X"0" & X"3e";
                    \$719_compbranch_arg\ := X"0000000" & X"4" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"88" =>
                    \$719_compbranch_id\ := X"0" & X"3f";
                    \$719_compbranch_arg\ := X"0000000" & X"5" & \$744_argument1\ & \$745_argument2\ & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when others =>
                    \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v1545\(0 to 15) & X"000" & X"3")));
                    state_var5312 <= pause_getI5292;
                  end case;
                when pause_getII5299 =>
                  \$744_argument1\ := \$code_value\;
                  \$v5297\ := eclat_resize(\$740\,8);
                  case \$v5297\ is
                  when X"0" & X"8" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & X"000" & X"1")));
                    state_var5312 <= pause_getI5170;
                  when X"12" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5174;
                  when X"13" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(16 to 47) & eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"14" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1") & eclat_resize(\$744_argument1\,16))));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5175;
                  when X"19" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(eclat_resize(\$744_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                    state_var5312 <= pause_getI5176;
                  when X"1e" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5180;
                  when X"1f" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(\$v1545\(96 to 103),31) & eclat_true;
                    state_var5312 <= pause_setI5183;
                  when X"20" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI5184;
                  when X"25" =>
                    \$711_apply_id\ := X"0" & X"27";
                    \$711_apply_arg\ := eclat_true & eclat_false & eclat_false & \$v1545\(96 to 103) & eclat_true & eclat_resize(\$744_argument1\,16) & X"000" & X"1" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"26" =>
                    \$711_apply_id\ := X"0" & X"28";
                    \$711_apply_arg\ := eclat_true & eclat_true & eclat_false & eclat_add(\$v1545\(96 to 103) & X"0" & X"1") & eclat_true & eclat_resize(\$744_argument1\,16) & X"000" & X"2" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"27" =>
                    \$711_apply_id\ := X"0" & X"29";
                    \$711_apply_arg\ := eclat_true & eclat_true & eclat_true & eclat_add(\$v1545\(96 to 103) & X"0" & X"2") & eclat_true & eclat_resize(\$744_argument1\,16) & X"000" & X"3" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"28" =>
                    \$v5194\ := eclat_gt(\$v1545\(96 to 103) & X"0" & X"0");
                    if \$v5194\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var5312 <= pause_getI5186;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16)) & X"000" & X"1")));
                      state_var5312 <= pause_getI5192;
                    end if;
                  when X"2a" =>
                    \$v5203\ := eclat_ge(\$v1545\(96 to 103) & eclat_resize(\$744_argument1\,8));
                    if \$v5203\(0) = '1' then
                      \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & eclat_sub(\$v1545\(96 to 103) & eclat_resize(\$744_argument1\,8)) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    else
                      \$710_id\ := X"0" & X"2b";
                      \$710_arg\ := \$v1545\(48 to 63) & \$v1545\(16 to 47) & \$v1545\(64 to 95) & X"f7" & eclat_resize(eclat_add(\$v1545\(96 to 103) & X"0" & X"3"),16) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                      state_var5312 <= \$710\;
                    end if;
                  when X"30" =>
                    \$712_offsetclosure_n_id\ := X"0" & X"2c";
                    \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16) & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    state_var5312 <= \$712_offsetclosure_n\;
                  when X"34" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5204;
                  when X"35" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$744_argument1\,16))));
                    state_var5312 <= pause_getI5205;
                  when X"36" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5209;
                  when X"39" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$744_argument1\,16))));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5210;
                  when X"3b" =>
                    \$716_make_block_n_id\ := X"0" & X"2e";
                    \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(48 to 63) & eclat_false & eclat_false & eclat_false & \$744_argument1\ & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$716_make_block_n\;
                  when X"3d" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5211;
                  when X"3f" =>
                    \$716_make_block_n_id\ := X"0" & X"30";
                    \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(48 to 63) & eclat_true & eclat_false & eclat_false & \$744_argument1\ & X"000" & X"1" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$716_make_block_n\;
                  when X"40" =>
                    \$716_make_block_n_id\ := X"0" & X"31";
                    \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(48 to 63) & eclat_true & eclat_true & eclat_false & \$744_argument1\ & X"000" & X"2" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$716_make_block_n\;
                  when X"41" =>
                    \$716_make_block_n_id\ := X"0" & X"32";
                    \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(48 to 63) & eclat_true & eclat_true & eclat_true & \$744_argument1\ & X"000" & X"3" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$716_make_block_n\;
                  when X"47" =>
                    eclat_skip(eclat_not(""&\$v1545\(47)));
                    
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & eclat_resize(\$744_argument1\,16)) & X"000" & X"1")));
                    state_var5312 <= pause_getI5212;
                  when X"4d" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5215;
                  when X"57" =>
                    \$v5221\ := ""&\$v1545\(47);
                    if \$v5221\(0) = '1' then
                      \$883_ofs\ := eclat_resize(\$v1545\(16 to 46),16);
                      \$code_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$883_ofs\)));
                      state_var5312 <= pause_getI5217;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v1545\(16 to 46),16)));
                      state_var5312 <= pause_getI5219;
                    end if;
                  when X"54" =>
                    \$v8\ := eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_resize(\$744_argument1\,16)) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"59" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(\$v1545\(96 to 103),31) & eclat_true;
                    state_var5312 <= pause_setI5225;
                  when X"5c" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(104 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"5d" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(64 to 95);
                    state_var5312 <= pause_setI5229;
                  when X"5e" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5234;
                  when X"5f" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5242;
                  when X"60" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5252;
                  when X"61" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5264;
                  when X"67" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$744_argument1\ & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"6c" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5266;
                  when X"7f" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(16 to 46) & \$744_argument1\) & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"80" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI5268;
                  when X"8b" =>
                    \$719_compbranch_id\ := X"0" & X"33";
                    \$719_compbranch_arg\ := X"0000000" & X"2" & \$744_argument1\ & \$v1545\(16 to 46) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when X"8c" =>
                    \$719_compbranch_id\ := X"0" & X"34";
                    \$719_compbranch_arg\ := X"0000000" & X"5" & \$744_argument1\ & \$v1545\(16 to 46) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_add(\$v1545\(0 to 15) & X"000" & X"3");
                    state_var5312 <= \$719_compbranch\;
                  when others =>
                    \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v1545\(0 to 15) & X"000" & X"2")));
                    state_var5312 <= pause_getI5295;
                  end case;
                when pause_getII5302 =>
                  \$740\ := \$code_value\;
                  \$v5300\ := eclat_resize(\$740\,8);
                  case \$v5300\ is
                  when X"0" & X"0" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI5049;
                  when X"0" & X"1" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                    state_var5312 <= pause_getI5051;
                  when X"0" & X"2" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"2") & X"000" & X"1")));
                    state_var5312 <= pause_getI5053;
                  when X"0" & X"3" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"3") & X"000" & X"1")));
                    state_var5312 <= pause_getI5055;
                  when X"0" & X"4" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"4") & X"000" & X"1")));
                    state_var5312 <= pause_getI5057;
                  when X"0" & X"5" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"5") & X"000" & X"1")));
                    state_var5312 <= pause_getI5059;
                  when X"0" & X"6" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"6") & X"000" & X"1")));
                    state_var5312 <= pause_getI5061;
                  when X"0" & X"7" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"7") & X"000" & X"1")));
                    state_var5312 <= pause_getI5063;
                  when X"0" & X"9" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5065;
                  when X"0" & X"a" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5066;
                  when X"0" & X"b" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5069;
                  when X"0" & X"c" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5072;
                  when X"0" & X"d" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5075;
                  when X"0" & X"e" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5078;
                  when X"0" & X"f" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5081;
                  when X"10" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5084;
                  when X"11" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5087;
                  when X"15" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                    state_var5312 <= pause_getI5088;
                  when X"16" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                    state_var5312 <= pause_getI5090;
                  when X"17" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                    state_var5312 <= pause_getI5092;
                  when X"18" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                    state_var5312 <= pause_getI5094;
                  when X"1a" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5098;
                  when X"1b" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5101;
                  when X"1c" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5104;
                  when X"1d" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5107;
                  when X"21" =>
                    \$711_apply_id\ := X"00" & X"c";
                    \$711_apply_arg\ := eclat_true & eclat_false & eclat_false & X"0" & X"0" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"22" =>
                    \$711_apply_id\ := X"00" & X"d";
                    \$711_apply_arg\ := eclat_true & eclat_true & eclat_false & X"0" & X"1" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"23" =>
                    \$711_apply_id\ := X"00" & X"e";
                    \$711_apply_arg\ := eclat_true & eclat_true & eclat_true & X"0" & X"2" & eclat_false & X"000" & X"0" & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(104 to 119);
                    state_var5312 <= \$711_apply\;
                  when X"29" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v1545\(64 to 94),16)));
                    state_var5312 <= pause_getI5110;
                  when X"2d" =>
                    \$712_offsetclosure_n_id\ := X"0" & X"10";
                    \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(48 to 63) & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    state_var5312 <= \$712_offsetclosure_n\;
                  when X"2e" =>
                    \$712_offsetclosure_n_id\ := X"0" & X"11";
                    \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(48 to 63) & X"000" & X"0" & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    state_var5312 <= \$712_offsetclosure_n\;
                  when X"2f" =>
                    \$712_offsetclosure_n_id\ := X"0" & X"12";
                    \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(48 to 63) & X"000" & X"2" & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    state_var5312 <= \$712_offsetclosure_n\;
                  when X"31" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5112;
                  when X"32" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5113;
                  when X"33" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5114;
                  when X"3a" =>
                    \$716_make_block_n_id\ := X"0" & X"16";
                    \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(48 to 63) & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                    state_var5312 <= \$716_make_block_n\;
                  when X"3c" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5115;
                  when X"43" =>
                    eclat_skip(eclat_not(""&\$v1545\(47)));
                    
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI5116;
                  when X"44" =>
                    eclat_skip(eclat_not(""&\$v1545\(47)));
                    
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"1") & X"000" & X"1")));
                    state_var5312 <= pause_getI5118;
                  when X"45" =>
                    eclat_skip(eclat_not(""&\$v1545\(47)));
                    
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"2") & X"000" & X"1")));
                    state_var5312 <= pause_getI5120;
                  when X"46" =>
                    eclat_skip(eclat_not(""&\$v1545\(47)));
                    
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(16 to 46),16) & X"000" & X"3") & X"000" & X"1")));
                    state_var5312 <= pause_getI5122;
                  when X"49" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5125;
                  when X"4a" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5128;
                  when X"4b" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5131;
                  when X"4c" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5134;
                  when X"4f" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$v1545\(16 to 46),16)));
                    state_var5312 <= pause_getI5136;
                  when X"50" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5140;
                  when X"51" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5145;
                  when X"52" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5149;
                  when X"53" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1")));
                    state_var5312 <= pause_getI5154;
                  when X"55" =>
                    \$717_branch_if_id\ := X"0" & X"18";
                    \$717_branch_if_arg\ := eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_add(\$v1545\(0 to 15) & X"000" & X"2");
                    state_var5312 <= \$717_branch_if\;
                  when X"56" =>
                    \$717_branch_if_id\ := X"0" & X"19";
                    \$717_branch_if_arg\ := eclat_true & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_add(\$v1545\(0 to 15) & X"000" & X"2");
                    state_var5312 <= \$717_branch_if\;
                  when X"58" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & 
                    eclat_if(eclat_eq(\$v1545\(16 to 46) & "000"& X"000000" & X"0") & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"5a" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$v1545\(48 to 63) & X"000" & X"1") & X"000" & X"1")));
                    state_var5312 <= pause_getI5156;
                  when X"5b" =>
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v1545\(104 to 119) & X"000" & X"1")));
                    state_var5312 <= pause_getI5164;
                  when X"63" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"64" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"65" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"66" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"68" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5166;
                  when X"69" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5167;
                  when X"6a" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5168;
                  when X"6b" =>
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v1545\(48 to 63)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v1545\(16 to 47);
                    state_var5312 <= pause_setI5169;
                  when X"6e" =>
                    \$713_binop_int_id\ := X"0" & X"1a";
                    \$713_binop_int_arg\ := X"0000000" & X"0" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"6f" =>
                    \$713_binop_int_id\ := X"0" & X"1b";
                    \$713_binop_int_arg\ := X"0000000" & X"1" & eclat_true & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"70" =>
                    \$713_binop_int_id\ := X"0" & X"1c";
                    \$713_binop_int_arg\ := X"0000000" & X"2" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"72" =>
                    \$713_binop_int_id\ := X"0" & X"1d";
                    \$713_binop_int_arg\ := X"0000000" & X"3" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"73" =>
                    \$713_binop_int_id\ := X"0" & X"1e";
                    \$713_binop_int_arg\ := X"0000000" & X"4" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"74" =>
                    \$713_binop_int_id\ := X"0" & X"1f";
                    \$713_binop_int_arg\ := X"0000000" & X"5" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"75" =>
                    \$713_binop_int_id\ := X"0" & X"20";
                    \$713_binop_int_arg\ := X"0000000" & X"6" & eclat_false & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$713_binop_int\;
                  when X"79" =>
                    \$715_binop_compare_id\ := X"0" & X"21";
                    \$715_binop_compare_arg\ := X"0000000" & X"0" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"7a" =>
                    \$715_binop_compare_id\ := X"0" & X"22";
                    \$715_binop_compare_arg\ := X"0000000" & X"1" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"7b" =>
                    \$715_binop_compare_id\ := X"0" & X"23";
                    \$715_binop_compare_arg\ := X"0000000" & X"2" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"7c" =>
                    \$715_binop_compare_id\ := X"0" & X"24";
                    \$715_binop_compare_arg\ := X"0000000" & X"3" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"7d" =>
                    \$715_binop_compare_id\ := X"0" & X"25";
                    \$715_binop_compare_arg\ := X"0000000" & X"4" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"7e" =>
                    \$715_binop_compare_id\ := X"0" & X"26";
                    \$715_binop_compare_arg\ := X"0000000" & X"5" & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121) & eclat_add(\$v1545\(0 to 15) & X"000" & X"1");
                    state_var5312 <= \$715_binop_compare\;
                  when X"81" =>
                    \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & 
                    eclat_if(""&\$v1545\(47) & "000"& X"000000" & X"1" & "000"& X"000000" & X"0") & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"8f" =>
                    eclat_print_string(of_string("STOP : "));
                    
                    \$v8\ := \$v1545\(0 to 15) & \$v1545\(16 to 47) & \$v1545\(48 to 63) & \$v1545\(64 to 119) & eclat_true & ""&\$v1545\(121);
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when others =>
                    \$code_ptr\ <= to_integer(unsigned(eclat_add(\$v1545\(0 to 15) & X"000" & X"1")));
                    state_var5312 <= pause_getI5298;
                  end case;
                when pause_setI5065 =>
                  \$ram_write_request\ <= '0';
                  \$v3660\ := eclat_unit;
                  \$1332_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(16 to 47) & \$1332_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5066 =>
                  \$ram_write_request\ <= '0';
                  \$v3661\ := eclat_unit;
                  \$5370_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$v1545\(16 to 47) & \$5370_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5069 =>
                  \$ram_write_request\ <= '0';
                  \$v3662\ := eclat_unit;
                  \$5372_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5372_sp\ & X"000" & X"1") & X"000" & X"1")));
                  state_var5312 <= pause_getI5067;
                when pause_setI5072 =>
                  \$ram_write_request\ <= '0';
                  \$v3663\ := eclat_unit;
                  \$5377_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5377_sp\ & X"000" & X"2") & X"000" & X"1")));
                  state_var5312 <= pause_getI5070;
                when pause_setI5075 =>
                  \$ram_write_request\ <= '0';
                  \$v3664\ := eclat_unit;
                  \$5382_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5382_sp\ & X"000" & X"3") & X"000" & X"1")));
                  state_var5312 <= pause_getI5073;
                when pause_setI5078 =>
                  \$ram_write_request\ <= '0';
                  \$v3665\ := eclat_unit;
                  \$5387_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5387_sp\ & X"000" & X"4") & X"000" & X"1")));
                  state_var5312 <= pause_getI5076;
                when pause_setI5081 =>
                  \$ram_write_request\ <= '0';
                  \$v3666\ := eclat_unit;
                  \$5392_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5392_sp\ & X"000" & X"5") & X"000" & X"1")));
                  state_var5312 <= pause_getI5079;
                when pause_setI5084 =>
                  \$ram_write_request\ <= '0';
                  \$v3667\ := eclat_unit;
                  \$5397_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5397_sp\ & X"000" & X"6") & X"000" & X"1")));
                  state_var5312 <= pause_getI5082;
                when pause_setI5087 =>
                  \$ram_write_request\ <= '0';
                  \$v3668\ := eclat_unit;
                  \$5402_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$5402_sp\ & X"000" & X"7") & X"000" & X"1")));
                  state_var5312 <= pause_getI5085;
                when pause_setI5098 =>
                  \$ram_write_request\ <= '0';
                  \$v3669\ := eclat_unit;
                  \$5427_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"1" & X"000" & X"1")) & X"000" & X"1")));
                  state_var5312 <= pause_getI5096;
                when pause_setI5101 =>
                  \$ram_write_request\ <= '0';
                  \$v3670\ := eclat_unit;
                  \$5434_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"2" & X"000" & X"1")) & X"000" & X"1")));
                  state_var5312 <= pause_getI5099;
                when pause_setI5104 =>
                  \$ram_write_request\ <= '0';
                  \$v3671\ := eclat_unit;
                  \$5441_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"3" & X"000" & X"1")) & X"000" & X"1")));
                  state_var5312 <= pause_getI5102;
                when pause_setI5107 =>
                  \$ram_write_request\ <= '0';
                  \$v3672\ := eclat_unit;
                  \$5448_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(X"000" & X"4" & X"000" & X"1")) & X"000" & X"1")));
                  state_var5312 <= pause_getI5105;
                when pause_setI5112 =>
                  \$ram_write_request\ <= '0';
                  \$v3673\ := eclat_unit;
                  \$5459_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$712_offsetclosure_n_id\ := X"0" & X"13";
                  \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5459_sp\ & eclat_sub(X"000" & X"0" & X"000" & X"2") & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  state_var5312 <= \$712_offsetclosure_n\;
                when pause_setI5113 =>
                  \$ram_write_request\ <= '0';
                  \$v3674\ := eclat_unit;
                  \$5461_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$712_offsetclosure_n_id\ := X"0" & X"14";
                  \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5461_sp\ & X"000" & X"0" & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  state_var5312 <= \$712_offsetclosure_n\;
                when pause_setI5114 =>
                  \$ram_write_request\ <= '0';
                  \$v3675\ := eclat_unit;
                  \$5463_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$712_offsetclosure_n_id\ := X"0" & X"15";
                  \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$5463_sp\ & X"000" & X"2" & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  state_var5312 <= \$712_offsetclosure_n\;
                when pause_setI5115 =>
                  \$ram_write_request\ <= '0';
                  \$v3676\ := eclat_unit;
                  \$975_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$716_make_block_n_id\ := X"0" & X"17";
                  \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & \$975_sp\ & eclat_false & eclat_false & eclat_false & "000"& X"000000" & X"0" & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                  state_var5312 <= \$716_make_block_n\;
                when pause_setI5124 =>
                  \$ram_write_request\ <= '0';
                  \$v3682\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3681\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5127 =>
                  \$ram_write_request\ <= '0';
                  \$v3684\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3683\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5130 =>
                  \$ram_write_request\ <= '0';
                  \$v3686\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3685\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5133 =>
                  \$ram_write_request\ <= '0';
                  \$v3688\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3687\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5142 =>
                  \$ram_write_request\ <= '0';
                  \$v3692\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3691\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5151 =>
                  \$ram_write_request\ <= '0';
                  \$v3696\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$v3695\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5166 =>
                  \$ram_write_request\ <= '0';
                  \$v3702\ := eclat_unit;
                  \$5557_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"0" & eclat_true & \$5557_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5167 =>
                  \$ram_write_request\ <= '0';
                  \$v3703\ := eclat_unit;
                  \$5560_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"1" & eclat_true & \$5560_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5168 =>
                  \$ram_write_request\ <= '0';
                  \$v3704\ := eclat_unit;
                  \$5563_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"2" & eclat_true & \$5563_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5169 =>
                  \$ram_write_request\ <= '0';
                  \$v3705\ := eclat_unit;
                  \$5566_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & "000"& X"000000" & X"3" & eclat_true & \$5566_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5174 =>
                  \$ram_write_request\ <= '0';
                  \$v3602\ := eclat_unit;
                  \$1312_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$1312_sp\ & eclat_resize(\$744_argument1\,16)) & X"000" & X"1")));
                  state_var5312 <= pause_getI5172;
                when pause_setI5175 =>
                  \$ram_write_request\ <= '0';
                  \$v3603\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5180 =>
                  \$ram_write_request\ <= '0';
                  \$v3604\ := eclat_unit;
                  \$1305_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v1545\(64 to 94),16) & eclat_sub(eclat_resize(\$744_argument1\,16) & X"000" & X"1")) & X"000" & X"1")));
                  state_var5312 <= pause_getI5178;
                when pause_setI5181 =>
                  \$ram_write_request\ <= '0';
                  \$v3605\ := eclat_unit;
                  \$820_sp\ := eclat_add(\$819_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(16 to 47) & \$820_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5182 =>
                  \$ram_write_request\ <= '0';
                  \$v3606\ := eclat_unit;
                  \$819_sp\ := eclat_add(\$814_sp\ & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$819_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_resize(\$744_argument1\,16)),31) & eclat_true;
                  state_var5312 <= pause_setI5181;
                when pause_setI5183 =>
                  \$ram_write_request\ <= '0';
                  \$v3607\ := eclat_unit;
                  \$814_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$814_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5182;
                when pause_setI5201 =>
                  \$ram_write_request\ <= '0';
                  \$v3613\ := eclat_unit;
                  \$720_w_id\ := X"0" & X"2a";
                  \$720_w_arg\ := X"0" & X"0" & \$v1545\(48 to 63) & \$v3611\(64 to 95) & \$v1545\(96 to 103);
                  state_var5312 <= \$720_w\;
                when pause_setI5202 =>
                  \$ram_write_request\ <= '0';
                  \$v3612\ := eclat_unit;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3611\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3611\(32 to 63);
                  state_var5312 <= pause_setI5201;
                when pause_setI5204 =>
                  \$ram_write_request\ <= '0';
                  \$v3617\ := eclat_unit;
                  \$1243_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$712_offsetclosure_n_id\ := X"0" & X"2d";
                  \$712_offsetclosure_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$1243_sp\ & eclat_resize(\$744_argument1\,16) & \$v1545\(64 to 95) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  state_var5312 <= \$712_offsetclosure_n\;
                when pause_setI5209 =>
                  \$ram_write_request\ <= '0';
                  \$v3618\ := eclat_unit;
                  \$875_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$744_argument1\,16))));
                  state_var5312 <= pause_getI5207;
                when pause_setI5210 =>
                  \$ram_write_request\ <= '0';
                  \$v3619\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5211 =>
                  \$ram_write_request\ <= '0';
                  \$v3620\ := eclat_unit;
                  \$879_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$716_make_block_n_id\ := X"0" & X"2f";
                  \$716_make_block_n_arg\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$879_sp\ & eclat_false & eclat_false & eclat_false & \$744_argument1\ & X"000" & X"0" & \$v1545\(16 to 47) & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$v1545\(120 to 121) & \$v1545\(104 to 119) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                  state_var5312 <= \$716_make_block_n\;
                when pause_setI5214 =>
                  \$ram_write_request\ <= '0';
                  \$v3623\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v3622\(32 to 47) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5222 =>
                  \$ram_write_request\ <= '0';
                  \$v3624\ := eclat_unit;
                  \$902_sp\ := eclat_add(\$901_sp\ & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$v1545\(16 to 47) & \$902_sp\ & \$v1545\(64 to 95) & \$v1545\(96 to 103) & \$902_sp\ & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5223 =>
                  \$ram_write_request\ <= '0';
                  \$v3625\ := eclat_unit;
                  \$901_sp\ := eclat_add(\$894_sp\ & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$901_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"1") & eclat_resize(\$744_argument1\,16)),31) & eclat_true;
                  state_var5312 <= pause_setI5222;
                when pause_setI5224 =>
                  \$ram_write_request\ <= '0';
                  \$v3626\ := eclat_unit;
                  \$894_sp\ := eclat_add(\$893_sp\ & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$894_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$v1545\(104 to 119),31) & eclat_true;
                  state_var5312 <= pause_setI5223;
                when pause_setI5225 =>
                  \$ram_write_request\ <= '0';
                  \$v3627\ := eclat_unit;
                  \$893_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$893_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v1545\(64 to 95);
                  state_var5312 <= pause_setI5224;
                when pause_setI5229 =>
                  \$ram_write_request\ <= '0';
                  \$v3631\ := eclat_unit;
                  \$903_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v5228\ := \$744_argument1\;
                  case \$v5228\ is
                  when others =>
                    eclat_print_string(of_string("unknown primitive"));
                    
                    \$v3628\ := "000"& X"000000" & X"1" & eclat_true & eclat_unit;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$903_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5226;
                  end case;
                when pause_setI5233 =>
                  \$ram_write_request\ <= '0';
                  \$v3636\ := eclat_unit;
                  \$912_sp\ := eclat_add(\$v3632\(32 to 47) & X"000" & X"1");
                  \$v5232\ := \$744_argument1\;
                  case \$v5232\ is
                  when others =>
                    eclat_print_string(of_string("unknown primitive"));
                    
                    \$v3633\ := "000"& X"000000" & X"1" & eclat_true & eclat_unit;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$912_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5230;
                  end case;
                when pause_setI5239 =>
                  \$ram_write_request\ <= '0';
                  \$v3642\ := eclat_unit;
                  \$923_sp\ := eclat_add(\$v3638\(32 to 47) & X"000" & X"1");
                  \$v5238\ := \$744_argument1\;
                  case \$v5238\ is
                  when others =>
                    eclat_print_string(of_string("unknown primitive"));
                    
                    \$v3639\ := "000"& X"000000" & X"1" & eclat_true & eclat_unit;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$923_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5236;
                  end case;
                when pause_setI5247 =>
                  \$ram_write_request\ <= '0';
                  \$v3649\ := eclat_unit;
                  \$936_sp\ := eclat_add(\$v3645\(32 to 47) & X"000" & X"1");
                  \$v5246\ := \$744_argument1\;
                  case \$v5246\ is
                  when others =>
                    eclat_print_string(of_string("unknown primitive"));
                    
                    \$v3646\ := "000"& X"000000" & X"1" & eclat_true & eclat_unit;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$936_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5244;
                  end case;
                when pause_setI5257 =>
                  \$ram_write_request\ <= '0';
                  \$v3657\ := eclat_unit;
                  \$951_sp\ := eclat_add(\$v3653\(32 to 47) & X"000" & X"1");
                  \$v5256\ := \$744_argument1\;
                  case \$v5256\ is
                  when others =>
                    eclat_print_string(of_string("unknown primitive"));
                    
                    \$v3654\ := "000"& X"000000" & X"1" & eclat_true & eclat_unit;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$951_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5254;
                  end case;
                when pause_setI5266 =>
                  \$ram_write_request\ <= '0';
                  \$v3658\ := eclat_unit;
                  \$1297_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & \$744_argument1\ & eclat_true & \$1297_sp\ & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5267 =>
                  \$ram_write_request\ <= '0';
                  \$v3659\ := eclat_unit;
                  \$v8\ := eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & "000"& X"000000" & X"1" & eclat_true & \$v1545\(48 to 63) & \$v1545\(64 to 119) & \$v1545\(120 to 121);
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5272 =>
                  \$ram_write_request\ <= '0';
                  \$v3597\ := eclat_unit;
                  \$v3595\ := \$v3596\(0 to 31) & \$v3596\(32 to 63) & \$v3596\(64 to 95);
                  \$722_fill_id\ := X"0" & X"36";
                  \$722_fill_arg\ := X"000" & X"1" & \$778_sp\ & eclat_resize(\$744_argument1\,16) & \$v3595\(64 to 95);
                  state_var5312 <= \$722_fill\;
                when pause_setI5273 =>
                  \$ram_write_request\ <= '0';
                  \$v3598\ := eclat_unit;
                  \$778_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$710_id\ := X"0" & X"37";
                  \$710_arg\ := \$778_sp\ & \$v1545\(16 to 47) & \$v1545\(64 to 95) & X"f7" & eclat_add(eclat_resize(\$744_argument1\,16) & X"000" & X"1") & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                  state_var5312 <= \$710\;
                when pause_setI5283 =>
                  \$ram_write_request\ <= '0';
                  \$v3599\ := eclat_unit;
                  \$792_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(X"3e80" & eclat_resize(\$744_argument1\,16))));
                  state_var5312 <= pause_getI5281;
                when pause_setI5284 =>
                  \$ram_write_request\ <= '0';
                  \$v3601\ := eclat_unit;
                  \$723_fill_id\ := X"0" & X"38";
                  \$723_fill_arg\ := X"000" & X"1" & \$v1545\(48 to 63) & eclat_resize(\$744_argument1\,16) & \$v3600\(64 to 95);
                  state_var5312 <= \$723_fill\;
                when pause_setI5285 =>
                  \$ram_write_request\ <= '0';
                  \$v3592\ := eclat_unit;
                  \$763_sp\ := eclat_add(\$762_sp\ & X"000" & X"1");
                  \$726_w3_id\ := X"0" & X"40";
                  \$726_w3_arg\ := X"000" & X"1" & \$763_sp\ & \$v3589\(64 to 95) & eclat_resize(\$744_argument1\,16);
                  state_var5312 <= \$726_w3\;
                when pause_setI5286 =>
                  \$ram_write_request\ <= '0';
                  \$v3590\ := eclat_unit;
                  \$724_w0_id\ := X"0" & X"42";
                  \$724_w0_arg\ := X"000" & X"0" & \$752_sp\ & eclat_resize(\$745_argument2\,16) & \$v3589\(64 to 95) & eclat_resize(\$744_argument1\,16);
                  state_var5312 <= \$724_w0\;
                when pause_setI5287 =>
                  \$ram_write_request\ <= '0';
                  \$v3593\ := eclat_unit;
                  \$752_sp\ := eclat_add(\$v1545\(48 to 63) & X"000" & X"1");
                  \$710_id\ := X"0" & X"43";
                  \$710_arg\ := \$752_sp\ & \$v1545\(16 to 47) & \$v1545\(64 to 95) & X"f7" & eclat_add(eclat_sub(eclat_mult(X"000" & X"2" & eclat_resize(\$744_argument1\,16)) & X"000" & X"1") & eclat_resize(\$745_argument2\,16)) & X"1770" & X"0" & X"fa0" & X"3e80" & X"0" & X"3e8";
                  state_var5312 <= \$710\;
                when pause_getI4922 =>
                  state_var5312 <= pause_getII4923;
                when pause_getII4923 =>
                  \$1636\ := \$ram_value\;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$706_loop_arg\(48 to 63) & \$706_loop_arg\(0 to 15))));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$1636\;
                  state_var5312 <= pause_setI4921;
                when pause_setI4921 =>
                  \$ram_write_request\ <= '0';
                  \$v3422\ := eclat_unit;
                  \$706_loop_arg\ := eclat_add(\$706_loop_arg\(0 to 15) & X"000" & X"1") & \$706_loop_arg\(16 to 31) & \$706_loop_arg\(32 to 47) & \$706_loop_arg\(48 to 63);
                  state_var5312 <= \$706_loop\;
                when pause_getI4929 =>
                  state_var5312 <= pause_getII4930;
                when pause_getI4932 =>
                  state_var5312 <= pause_getII4933;
                when pause_getI4935 =>
                  state_var5312 <= pause_getII4936;
                when pause_getII4930 =>
                  \$1618_hd\ := \$ram_value\;
                  \$1620\ := eclat_resize(eclat_lsr(\$1618_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                  eclat_print_string(of_string("bloc "));
                  
                  eclat_print_int(eclat_resize(\$1603\(0 to 30),16));
                  
                  eclat_print_string(of_string(" of size "));
                  
                  eclat_print_int(eclat_add(\$1620\ & X"000" & X"1"));
                  
                  eclat_print_string(of_string(" from "));
                  
                  eclat_print_int(eclat_resize(\$1603\(0 to 30),16));
                  
                  eclat_print_string(of_string(" to "));
                  
                  eclat_print_int(\$707_copy_root_in_ram_arg\(32 to 47));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$ram_ptr_write\ <= to_integer(unsigned(\$707_copy_root_in_ram_arg\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$1618_hd\;
                  state_var5312 <= pause_setI4928;
                when pause_getII4933 =>
                  \$1616_w\ := \$ram_value\;
                  \$v4931\ := eclat_if(eclat_not(""&\$1616_w\(31)) & 
                              eclat_if(eclat_le(\$707_copy_root_in_ram_arg\(64 to 79) & eclat_resize(\$1616_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$1616_w\(0 to 30),16) & eclat_add(\$707_copy_root_in_ram_arg\(64 to 79) & \$707_copy_root_in_ram_arg\(80 to 95))) & eclat_false) & eclat_false);
                  if \$v4931\(0) = '1' then
                    \$v3427\ := \$1616_w\ & \$707_copy_root_in_ram_arg\(32 to 47);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$707_copy_root_in_ram_arg\(0 to 15)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3427\(0 to 31);
                    state_var5312 <= pause_setI4925;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$1603\(0 to 30),16)));
                    state_var5312 <= pause_getI4929;
                  end if;
                when pause_getII4936 =>
                  \$1603\ := \$ram_value\;
                  \$v4934\ := eclat_not(eclat_if(eclat_not(""&\$1603\(31)) & 
                                        eclat_if(eclat_le(\$707_copy_root_in_ram_arg\(48 to 63) & eclat_resize(\$1603\(0 to 30),16)) & eclat_lt(eclat_resize(\$1603\(0 to 30),16) & eclat_add(\$707_copy_root_in_ram_arg\(48 to 63) & \$707_copy_root_in_ram_arg\(80 to 95))) & eclat_false) & eclat_false));
                  if \$v4934\(0) = '1' then
                    \$v3427\ := \$1603\ & \$707_copy_root_in_ram_arg\(32 to 47);
                    \$ram_ptr_write\ <= to_integer(unsigned(\$707_copy_root_in_ram_arg\(0 to 15)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3427\(0 to 31);
                    state_var5312 <= pause_setI4925;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$1603\(0 to 30),16) & X"000" & X"1")));
                    state_var5312 <= pause_getI4932;
                  end if;
                when pause_setI4925 =>
                  \$ram_write_request\ <= '0';
                  \$v3428\ := eclat_unit;
                  eclat_print_string(of_string(" next="));
                  
                  eclat_print_int(\$v3427\(32 to 47));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$707_copy_root_in_ram_arg\ := eclat_add(\$707_copy_root_in_ram_arg\(0 to 15) & X"000" & X"1") & \$707_copy_root_in_ram_arg\(16 to 31) & \$v3427\(32 to 47) & \$707_copy_root_in_ram_arg\(48 to 63) & \$707_copy_root_in_ram_arg\(64 to 79) & \$707_copy_root_in_ram_arg\(80 to 95);
                  state_var5312 <= \$707_copy_root_in_ram\;
                when pause_setI4926 =>
                  \$ram_write_request\ <= '0';
                  \$v3444\ := eclat_unit;
                  \$v3427\ := eclat_resize(\$707_copy_root_in_ram_arg\(32 to 47),31) & eclat_false & eclat_add(\$707_copy_root_in_ram_arg\(32 to 47) & eclat_add(\$1620\ & X"000" & X"1"));
                  \$ram_ptr_write\ <= to_integer(unsigned(\$707_copy_root_in_ram_arg\(0 to 15)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3427\(0 to 31);
                  state_var5312 <= pause_setI4925;
                when pause_setI4927 =>
                  \$ram_write_request\ <= '0';
                  \$v3443\ := eclat_unit;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$1603\(0 to 30),16) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$707_copy_root_in_ram_arg\(32 to 47),31) & eclat_false;
                  state_var5312 <= pause_setI4926;
                when pause_setI4928 =>
                  \$ram_write_request\ <= '0';
                  \$v3441\ := eclat_unit;
                  \$706_loop_id\ := X"00" & X"1";
                  \$706_loop_arg\ := X"000" & X"1" & eclat_resize(\$1603\(0 to 30),16) & eclat_add(\$1620\ & X"000" & X"1") & \$707_copy_root_in_ram_arg\(32 to 47);
                  state_var5312 <= \$706_loop\;
                when pause_getI4942 =>
                  state_var5312 <= pause_getII4943;
                when pause_getI4945 =>
                  state_var5312 <= pause_getII4946;
                when pause_getI4948 =>
                  state_var5312 <= pause_getII4949;
                when pause_getII4943 =>
                  \$5083_hd\ := \$ram_value\;
                  \$5085\ := eclat_resize(eclat_lsr(\$5083_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                  eclat_print_string(of_string("bloc "));
                  
                  eclat_print_int(eclat_resize(\$1592\(0 to 30),16));
                  
                  eclat_print_string(of_string(" of size "));
                  
                  eclat_print_int(eclat_add(\$5085\ & X"000" & X"1"));
                  
                  eclat_print_string(of_string(" from "));
                  
                  eclat_print_int(eclat_resize(\$1592\(0 to 30),16));
                  
                  eclat_print_string(of_string(" to "));
                  
                  eclat_print_int(\$708_loop_arg\(16 to 31));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$ram_ptr_write\ <= to_integer(unsigned(\$708_loop_arg\(16 to 31)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$5083_hd\;
                  state_var5312 <= pause_setI4941;
                when pause_getII4946 =>
                  \$5081_w\ := \$ram_value\;
                  \$v4944\ := eclat_if(eclat_not(""&\$5081_w\(31)) & 
                              eclat_if(eclat_le(\$708_loop_arg\(64 to 79) & eclat_resize(\$5081_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$5081_w\(0 to 30),16) & eclat_add(\$708_loop_arg\(64 to 79) & \$708_loop_arg\(96 to 111))) & eclat_false) & eclat_false);
                  if \$v4944\(0) = '1' then
                    \$v3446\ := \$5081_w\ & \$708_loop_arg\(16 to 31);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$708_loop_arg\(80 to 95) & \$708_loop_arg\(0 to 15))));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3446\(0 to 31);
                    state_var5312 <= pause_setI4938;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$1592\(0 to 30),16)));
                    state_var5312 <= pause_getI4942;
                  end if;
                when pause_getII4949 =>
                  \$1592\ := \$ram_value\;
                  \$v4947\ := eclat_not(eclat_if(eclat_not(""&\$1592\(31)) & 
                                        eclat_if(eclat_le(\$708_loop_arg\(48 to 63) & eclat_resize(\$1592\(0 to 30),16)) & eclat_lt(eclat_resize(\$1592\(0 to 30),16) & eclat_add(\$708_loop_arg\(48 to 63) & \$708_loop_arg\(96 to 111))) & eclat_false) & eclat_false));
                  if \$v4947\(0) = '1' then
                    \$v3446\ := \$1592\ & \$708_loop_arg\(16 to 31);
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$708_loop_arg\(80 to 95) & \$708_loop_arg\(0 to 15))));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3446\(0 to 31);
                    state_var5312 <= pause_setI4938;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$1592\(0 to 30),16) & X"000" & X"1")));
                    state_var5312 <= pause_getI4945;
                  end if;
                when pause_setI4938 =>
                  \$ram_write_request\ <= '0';
                  \$v3447\ := eclat_unit;
                  \$708_loop_arg\ := eclat_add(\$708_loop_arg\(0 to 15) & X"000" & X"1") & \$v3446\(32 to 47) & \$708_loop_arg\(32 to 47) & \$708_loop_arg\(48 to 63) & \$708_loop_arg\(64 to 79) & \$708_loop_arg\(80 to 95) & \$708_loop_arg\(96 to 111);
                  state_var5312 <= \$708_loop\;
                when pause_setI4939 =>
                  \$ram_write_request\ <= '0';
                  \$v3460\ := eclat_unit;
                  \$v3446\ := eclat_resize(\$708_loop_arg\(16 to 31),31) & eclat_false & eclat_add(\$708_loop_arg\(16 to 31) & eclat_add(\$5085\ & X"000" & X"1"));
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(\$708_loop_arg\(80 to 95) & \$708_loop_arg\(0 to 15))));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3446\(0 to 31);
                  state_var5312 <= pause_setI4938;
                when pause_setI4940 =>
                  \$ram_write_request\ <= '0';
                  \$v3459\ := eclat_unit;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$1592\(0 to 30),16) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$708_loop_arg\(16 to 31),31) & eclat_false;
                  state_var5312 <= pause_setI4939;
                when pause_setI4941 =>
                  \$ram_write_request\ <= '0';
                  \$v3457\ := eclat_unit;
                  \$706_loop_id\ := X"00" & X"2";
                  \$706_loop_arg\ := X"000" & X"1" & eclat_resize(\$1592\(0 to 30),16) & eclat_add(\$5085\ & X"000" & X"1") & \$708_loop_arg\(16 to 31);
                  state_var5312 <= \$706_loop\;
                when pause_getI4951 =>
                  state_var5312 <= pause_getII4952;
                when pause_getII4952 =>
                  \$1576\ := \$ram_value\;
                  \$1579\ := eclat_resize(eclat_lsr(eclat_resize(eclat_resize(\$1576\(0 to 30),16),31) & "000"& X"000000" & X"2"),16);
                  \$708_loop_id\ := X"00" & X"3";
                  \$708_loop_arg\ := X"000" & X"1" & \$709_aux_arg\(16 to 31) & eclat_add(\$1579\ & X"000" & X"1") & \$709_aux_arg\(32 to 47) & \$709_aux_arg\(48 to 63) & \$709_aux_arg\(0 to 15) & \$709_aux_arg\(64 to 79);
                  state_var5312 <= \$708_loop\;
                when pause_getI4955 =>
                  state_var5312 <= pause_getII4956;
                when pause_getI4960 =>
                  state_var5312 <= pause_getII4961;
                when pause_getI4963 =>
                  state_var5312 <= pause_getII4964;
                when pause_getI4969 =>
                  state_var5312 <= pause_getII4970;
                when pause_getI4972 =>
                  state_var5312 <= pause_getII4973;
                when pause_getII4956 =>
                  \$1566\ := \$global_end_value\;
                  \$707_copy_root_in_ram_id\ := X"00" & X"5";
                  \$707_copy_root_in_ram_arg\ := \$710_arg\(136 to 151) & \$1566\ & \$1565_next\ & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                  state_var5312 <= \$707_copy_root_in_ram\;
                when pause_getII4961 =>
                  \$5112_hd\ := \$ram_value\;
                  \$5114\ := eclat_resize(eclat_lsr(\$5112_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                  eclat_print_string(of_string("bloc "));
                  
                  eclat_print_int(eclat_resize(\$710_arg\(48 to 78),16));
                  
                  eclat_print_string(of_string(" of size "));
                  
                  eclat_print_int(eclat_add(\$5114\ & X"000" & X"1"));
                  
                  eclat_print_string(of_string(" from "));
                  
                  eclat_print_int(eclat_resize(\$710_arg\(48 to 78),16));
                  
                  eclat_print_string(of_string(" to "));
                  
                  eclat_print_int(\$v3486\(32 to 47));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3486\(32 to 47)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$5112_hd\;
                  state_var5312 <= pause_setI4959;
                when pause_getII4964 =>
                  \$5110_w\ := \$ram_value\;
                  \$v4962\ := eclat_if(eclat_not(""&\$5110_w\(31)) & 
                              eclat_if(eclat_le(\$v3419\(112 to 127) & eclat_resize(\$5110_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$5110_w\(0 to 30),16) & eclat_add(\$v3419\(112 to 127) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false);
                  if \$v4962\(0) = '1' then
                    \$v3487\ := \$5110_w\ & \$v3486\(32 to 47);
                    \$707_copy_root_in_ram_id\ := X"00" & X"6";
                    \$707_copy_root_in_ram_arg\ := \$710_arg\(152 to 167) & \$710_arg\(0 to 15) & \$v3487\(32 to 47) & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                    state_var5312 <= \$707_copy_root_in_ram\;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$710_arg\(48 to 78),16)));
                    state_var5312 <= pause_getI4960;
                  end if;
                when pause_getII4970 =>
                  \$5139_hd\ := \$ram_value\;
                  \$5141\ := eclat_resize(eclat_lsr(\$5139_hd\(0 to 30) & "000"& X"000000" & X"2"),16);
                  eclat_print_string(of_string("bloc "));
                  
                  eclat_print_int(eclat_resize(\$710_arg\(16 to 46),16));
                  
                  eclat_print_string(of_string(" of size "));
                  
                  eclat_print_int(eclat_add(\$5141\ & X"000" & X"1"));
                  
                  eclat_print_string(of_string(" from "));
                  
                  eclat_print_int(eclat_resize(\$710_arg\(16 to 46),16));
                  
                  eclat_print_string(of_string(" to "));
                  
                  eclat_print_int(\$v3419\(112 to 127));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$ram_ptr_write\ <= to_integer(unsigned(\$v3419\(112 to 127)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$5139_hd\;
                  state_var5312 <= pause_setI4968;
                when pause_getII4973 =>
                  \$5137_w\ := \$ram_value\;
                  \$v4971\ := eclat_if(eclat_not(""&\$5137_w\(31)) & 
                              eclat_if(eclat_le(\$v3419\(112 to 127) & eclat_resize(\$5137_w\(0 to 30),16)) & eclat_lt(eclat_resize(\$5137_w\(0 to 30),16) & eclat_add(\$v3419\(112 to 127) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false);
                  if \$v4971\(0) = '1' then
                    \$v3486\ := \$5137_w\ & \$v3419\(112 to 127);
                    \$v4965\ := eclat_not(eclat_if(eclat_not(""&\$710_arg\(79)) & 
                                          eclat_if(eclat_le(\$v3419\(96 to 111) & eclat_resize(\$710_arg\(48 to 78),16)) & eclat_lt(eclat_resize(\$710_arg\(48 to 78),16) & eclat_add(\$v3419\(96 to 111) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false));
                    if \$v4965\(0) = '1' then
                      \$v3487\ := \$710_arg\(48 to 79) & \$v3486\(32 to 47);
                      \$707_copy_root_in_ram_id\ := X"00" & X"6";
                      \$707_copy_root_in_ram_arg\ := \$710_arg\(152 to 167) & \$710_arg\(0 to 15) & \$v3487\(32 to 47) & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                      state_var5312 <= \$707_copy_root_in_ram\;
                    else
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(48 to 78),16) & X"000" & X"1")));
                      state_var5312 <= pause_getI4963;
                    end if;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_resize(\$710_arg\(16 to 46),16)));
                    state_var5312 <= pause_getI4969;
                  end if;
                when pause_setI4954 =>
                  \$ram_write_request\ <= '0';
                  \$v3472\ := eclat_unit;
                  \$710_result\ := \$v3468\(0 to 31) & \$v3468\(32 to 63) & eclat_resize(\$v3468\(64 to 79),31) & eclat_false;
                  case \$710_id\ is
                  when X"00" & X"a" =>
                    \$v3547\ := \$710_result\;
                    \$v5014\ := ""&\$716_make_block_n_arg\(32);
                    if \$v5014\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3547\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v3547\(0 to 31);
                      state_var5312 <= pause_setI5013;
                    else
                      \$v3548\ := eclat_unit;
                      \$v5012\ := ""&\$716_make_block_n_arg\(33);
                      if \$v5012\(0) = '1' then
                        \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$716_make_block_n_arg\(16 to 31) & X"000" & X"1")));
                        state_var5312 <= pause_getI5010;
                      else
                        \$1179_sp\ := \$716_make_block_n_arg\(16 to 31);
                        \$v5008\ := ""&\$716_make_block_n_arg\(34);
                        if \$v5008\(0) = '1' then
                          \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$1179_sp\ & X"000" & X"1")));
                          state_var5312 <= pause_getI5006;
                        else
                          \$1180_sp\ := \$1179_sp\;
                          \$716_make_block_n_result\ := \$716_make_block_n_arg\(0 to 15) & \$v3547\(64 to 95) & \$1180_sp\ & \$v3547\(32 to 63) & \$716_make_block_n_arg\(146 to 153) & \$716_make_block_n_arg\(156 to 171) & \$716_make_block_n_arg\(154 to 155);
                          \$v8\ := \$716_make_block_n_result\;
                          \$v1549\ := \$v8\ & eclat_true;
                          result4918 := eclat_unit;
                          rdy4919 := eclat_true;
                          state_var5312 <= compute4920;
                        end if;
                      end if;
                    end if;
                  when X"0" & X"2b" =>
                    \$v3611\ := \$710_result\;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3611\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_sub(eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & X"000" & X"3"),31) & eclat_true;
                    state_var5312 <= pause_setI5202;
                  when X"0" & X"37" =>
                    \$v3596\ := \$710_result\;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3596\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"2") & eclat_resize(\$745_argument2\,16)),31) & eclat_true;
                    state_var5312 <= pause_setI5272;
                  when X"0" & X"39" =>
                    \$v3600\ := \$710_result\;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3600\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3600\(0 to 31);
                    state_var5312 <= pause_setI5284;
                  when X"0" & X"43" =>
                    \$v3589\ := \$710_result\;
                    \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3589\(64 to 94),16) & X"000" & X"0") & X"000" & X"1")));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(eclat_add(eclat_add(\$v1545\(0 to 15) & X"000" & X"3") & eclat_resize(\$746_argument3\,16)),31) & eclat_true;
                    state_var5312 <= pause_setI5286;
                  when others =>
                    
                  end case;
                when pause_setI4957 =>
                  \$ram_write_request\ <= '0';
                  \$v3506\ := eclat_unit;
                  \$v3487\ := eclat_resize(\$v3486\(32 to 47),31) & eclat_false & eclat_add(\$v3486\(32 to 47) & eclat_add(\$5114\ & X"000" & X"1"));
                  \$707_copy_root_in_ram_id\ := X"00" & X"6";
                  \$707_copy_root_in_ram_arg\ := \$710_arg\(152 to 167) & \$710_arg\(0 to 15) & \$v3487\(32 to 47) & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                  state_var5312 <= \$707_copy_root_in_ram\;
                when pause_setI4958 =>
                  \$ram_write_request\ <= '0';
                  \$v3505\ := eclat_unit;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(48 to 78),16) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$v3486\(32 to 47),31) & eclat_false;
                  state_var5312 <= pause_setI4957;
                when pause_setI4959 =>
                  \$ram_write_request\ <= '0';
                  \$v3503\ := eclat_unit;
                  \$706_loop_id\ := X"00" & X"7";
                  \$706_loop_arg\ := X"000" & X"1" & eclat_resize(\$710_arg\(48 to 78),16) & eclat_add(\$5114\ & X"000" & X"1") & \$v3486\(32 to 47);
                  state_var5312 <= \$706_loop\;
                when pause_setI4966 =>
                  \$ram_write_request\ <= '0';
                  \$v3519\ := eclat_unit;
                  \$v3486\ := eclat_resize(\$v3419\(112 to 127),31) & eclat_false & eclat_add(\$v3419\(112 to 127) & eclat_add(\$5141\ & X"000" & X"1"));
                  \$v4965\ := eclat_not(eclat_if(eclat_not(""&\$710_arg\(79)) & 
                                        eclat_if(eclat_le(\$v3419\(96 to 111) & eclat_resize(\$710_arg\(48 to 78),16)) & eclat_lt(eclat_resize(\$710_arg\(48 to 78),16) & eclat_add(\$v3419\(96 to 111) & \$710_arg\(104 to 119))) & eclat_false) & eclat_false));
                  if \$v4965\(0) = '1' then
                    \$v3487\ := \$710_arg\(48 to 79) & \$v3486\(32 to 47);
                    \$707_copy_root_in_ram_id\ := X"00" & X"6";
                    \$707_copy_root_in_ram_arg\ := \$710_arg\(152 to 167) & \$710_arg\(0 to 15) & \$v3487\(32 to 47) & \$v3419\(96 to 111) & \$v3419\(112 to 127) & \$710_arg\(104 to 119);
                    state_var5312 <= \$707_copy_root_in_ram\;
                  else
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(48 to 78),16) & X"000" & X"1")));
                    state_var5312 <= pause_getI4963;
                  end if;
                when pause_setI4967 =>
                  \$ram_write_request\ <= '0';
                  \$v3518\ := eclat_unit;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_resize(\$710_arg\(16 to 46),16) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$v3419\(112 to 127),31) & eclat_false;
                  state_var5312 <= pause_setI4966;
                when pause_setI4968 =>
                  \$ram_write_request\ <= '0';
                  \$v3516\ := eclat_unit;
                  \$706_loop_id\ := X"00" & X"8";
                  \$706_loop_arg\ := X"000" & X"1" & eclat_resize(\$710_arg\(16 to 46),16) & eclat_add(\$5141\ & X"000" & X"1") & \$v3419\(112 to 127);
                  state_var5312 <= \$706_loop\;
                when pause_getI4977 =>
                  state_var5312 <= pause_getII4978;
                when pause_getI4989 =>
                  state_var5312 <= pause_getII4990;
                when pause_getI4992 =>
                  state_var5312 <= pause_getII4993;
                when pause_getI4995 =>
                  state_var5312 <= pause_getII4996;
                when pause_getII4978 =>
                  \$1279\ := \$ram_value\;
                  \$711_apply_result\ := eclat_resize(\$1279\(0 to 30),16) & \$711_apply_arg\(44 to 75) & \$1278_sp\ & \$711_apply_arg\(44 to 75) & \$711_apply_arg\(3 to 10) & \$711_apply_arg\(150 to 165) & \$711_apply_arg\(132 to 133);
                  \$v8\ := \$711_apply_result\;
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getII4990 =>
                  \$1822_v\ := \$ram_value\;
                  \$v3530\ := \$1822_v\ & eclat_sub(\$v3529\(32 to 47) & X"000" & X"1");
                  \$v4988\ := ""&\$711_apply_arg\(11);
                  if \$v4988\(0) = '1' then
                    \$1275_sp\ := eclat_add(eclat_sub(\$v3530\(32 to 47) & \$711_apply_arg\(12 to 27)) & \$711_apply_arg\(28 to 43));
                    \$v4984\ := ""&\$711_apply_arg\(2);
                    if \$v4984\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v3530\(0 to 31);
                      state_var5312 <= pause_setI4983;
                    else
                      \$1276_sp\ := \$1275_sp\;
                      \$v4982\ := ""&\$711_apply_arg\(1);
                      if \$v4982\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v3529\(0 to 31);
                        state_var5312 <= pause_setI4981;
                      else
                        \$1277_sp\ := \$1276_sp\;
                        \$v4980\ := ""&\$711_apply_arg\(0);
                        if \$v4980\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v3528\(0 to 31);
                          state_var5312 <= pause_setI4979;
                        else
                          \$1278_sp\ := \$1277_sp\;
                          \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                          state_var5312 <= pause_getI4977;
                        end if;
                      end if;
                    end if;
                  else
                    \$ram_ptr_write\ <= to_integer(unsigned(\$v3530\(32 to 47)));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= eclat_resize(\$711_apply_arg\(124 to 131),31) & eclat_true;
                    state_var5312 <= pause_setI4987;
                  end if;
                when pause_getII4993 =>
                  \$5166_v\ := \$ram_value\;
                  \$v3529\ := \$5166_v\ & eclat_sub(\$v3528\(32 to 47) & X"000" & X"1");
                  \$v4991\ := ""&\$711_apply_arg\(2);
                  if \$v4991\(0) = '1' then
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3529\(32 to 47) & X"000" & X"1")));
                    state_var5312 <= pause_getI4989;
                  else
                    \$v3530\ := "000"& X"000000" & X"1" & eclat_true & \$v3529\(32 to 47);
                    \$v4988\ := ""&\$711_apply_arg\(11);
                    if \$v4988\(0) = '1' then
                      \$1275_sp\ := eclat_add(eclat_sub(\$v3530\(32 to 47) & \$711_apply_arg\(12 to 27)) & \$711_apply_arg\(28 to 43));
                      \$v4984\ := ""&\$711_apply_arg\(2);
                      if \$v4984\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v3530\(0 to 31);
                        state_var5312 <= pause_setI4983;
                      else
                        \$1276_sp\ := \$1275_sp\;
                        \$v4982\ := ""&\$711_apply_arg\(1);
                        if \$v4982\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v3529\(0 to 31);
                          state_var5312 <= pause_setI4981;
                        else
                          \$1277_sp\ := \$1276_sp\;
                          \$v4980\ := ""&\$711_apply_arg\(0);
                          if \$v4980\(0) = '1' then
                            \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$v3528\(0 to 31);
                            state_var5312 <= pause_setI4979;
                          else
                            \$1278_sp\ := \$1277_sp\;
                            \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                            state_var5312 <= pause_getI4977;
                          end if;
                        end if;
                      end if;
                    else
                      \$ram_ptr_write\ <= to_integer(unsigned(\$v3530\(32 to 47)));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= eclat_resize(\$711_apply_arg\(124 to 131),31) & eclat_true;
                      state_var5312 <= pause_setI4987;
                    end if;
                  end if;
                when pause_getII4996 =>
                  \$5168_v\ := \$ram_value\;
                  \$v3528\ := \$5168_v\ & eclat_sub(\$711_apply_arg\(76 to 91) & X"000" & X"1");
                  \$v4994\ := ""&\$711_apply_arg\(1);
                  if \$v4994\(0) = '1' then
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3528\(32 to 47) & X"000" & X"1")));
                    state_var5312 <= pause_getI4992;
                  else
                    \$v3529\ := "000"& X"000000" & X"1" & eclat_true & \$v3528\(32 to 47);
                    \$v4991\ := ""&\$711_apply_arg\(2);
                    if \$v4991\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$v3529\(32 to 47) & X"000" & X"1")));
                      state_var5312 <= pause_getI4989;
                    else
                      \$v3530\ := "000"& X"000000" & X"1" & eclat_true & \$v3529\(32 to 47);
                      \$v4988\ := ""&\$711_apply_arg\(11);
                      if \$v4988\(0) = '1' then
                        \$1275_sp\ := eclat_add(eclat_sub(\$v3530\(32 to 47) & \$711_apply_arg\(12 to 27)) & \$711_apply_arg\(28 to 43));
                        \$v4984\ := ""&\$711_apply_arg\(2);
                        if \$v4984\(0) = '1' then
                          \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                          \$ram_write_request\ <= '1';
                          \$ram_write\ <= \$v3530\(0 to 31);
                          state_var5312 <= pause_setI4983;
                        else
                          \$1276_sp\ := \$1275_sp\;
                          \$v4982\ := ""&\$711_apply_arg\(1);
                          if \$v4982\(0) = '1' then
                            \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                            \$ram_write_request\ <= '1';
                            \$ram_write\ <= \$v3529\(0 to 31);
                            state_var5312 <= pause_setI4981;
                          else
                            \$1277_sp\ := \$1276_sp\;
                            \$v4980\ := ""&\$711_apply_arg\(0);
                            if \$v4980\(0) = '1' then
                              \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                              \$ram_write_request\ <= '1';
                              \$ram_write\ <= \$v3528\(0 to 31);
                              state_var5312 <= pause_setI4979;
                            else
                              \$1278_sp\ := \$1277_sp\;
                              \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                              state_var5312 <= pause_getI4977;
                            end if;
                          end if;
                        end if;
                      else
                        \$ram_ptr_write\ <= to_integer(unsigned(\$v3530\(32 to 47)));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= eclat_resize(\$711_apply_arg\(124 to 131),31) & eclat_true;
                        state_var5312 <= pause_setI4987;
                      end if;
                    end if;
                  end if;
                when pause_setI4979 =>
                  \$ram_write_request\ <= '0';
                  \$v3531\ := eclat_unit;
                  \$1278_sp\ := eclat_add(\$1277_sp\ & X"000" & X"1");
                  \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                  state_var5312 <= pause_getI4977;
                when pause_setI4981 =>
                  \$ram_write_request\ <= '0';
                  \$v3532\ := eclat_unit;
                  \$1277_sp\ := eclat_add(\$1276_sp\ & X"000" & X"1");
                  \$v4980\ := ""&\$711_apply_arg\(0);
                  if \$v4980\(0) = '1' then
                    \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3528\(0 to 31);
                    state_var5312 <= pause_setI4979;
                  else
                    \$1278_sp\ := \$1277_sp\;
                    \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                    state_var5312 <= pause_getI4977;
                  end if;
                when pause_setI4983 =>
                  \$ram_write_request\ <= '0';
                  \$v3533\ := eclat_unit;
                  \$1276_sp\ := eclat_add(\$1275_sp\ & X"000" & X"1");
                  \$v4982\ := ""&\$711_apply_arg\(1);
                  if \$v4982\(0) = '1' then
                    \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3529\(0 to 31);
                    state_var5312 <= pause_setI4981;
                  else
                    \$1277_sp\ := \$1276_sp\;
                    \$v4980\ := ""&\$711_apply_arg\(0);
                    if \$v4980\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v3528\(0 to 31);
                      state_var5312 <= pause_setI4979;
                    else
                      \$1278_sp\ := \$1277_sp\;
                      \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                      state_var5312 <= pause_getI4977;
                    end if;
                  end if;
                when pause_setI4985 =>
                  \$ram_write_request\ <= '0';
                  \$v3534\ := eclat_unit;
                  \$1288_sp\ := eclat_add(\$1285_sp\ & X"000" & X"1");
                  \$1275_sp\ := \$1288_sp\;
                  \$v4984\ := ""&\$711_apply_arg\(2);
                  if \$v4984\(0) = '1' then
                    \$ram_ptr_write\ <= to_integer(unsigned(\$1275_sp\));
                    \$ram_write_request\ <= '1';
                    \$ram_write\ <= \$v3530\(0 to 31);
                    state_var5312 <= pause_setI4983;
                  else
                    \$1276_sp\ := \$1275_sp\;
                    \$v4982\ := ""&\$711_apply_arg\(1);
                    if \$v4982\(0) = '1' then
                      \$ram_ptr_write\ <= to_integer(unsigned(\$1276_sp\));
                      \$ram_write_request\ <= '1';
                      \$ram_write\ <= \$v3529\(0 to 31);
                      state_var5312 <= pause_setI4981;
                    else
                      \$1277_sp\ := \$1276_sp\;
                      \$v4980\ := ""&\$711_apply_arg\(0);
                      if \$v4980\(0) = '1' then
                        \$ram_ptr_write\ <= to_integer(unsigned(\$1277_sp\));
                        \$ram_write_request\ <= '1';
                        \$ram_write\ <= \$v3528\(0 to 31);
                        state_var5312 <= pause_setI4979;
                      else
                        \$1278_sp\ := \$1277_sp\;
                        \$ram_ptr\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$711_apply_arg\(44 to 74),16) & X"000" & X"0") & X"000" & X"1")));
                        state_var5312 <= pause_getI4977;
                      end if;
                    end if;
                  end if;
                when pause_setI4986 =>
                  \$ram_write_request\ <= '0';
                  \$v3535\ := eclat_unit;
                  \$1285_sp\ := eclat_add(\$1284_sp\ & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$1285_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= eclat_resize(\$711_apply_arg\(134 to 149),31) & eclat_true;
                  state_var5312 <= pause_setI4985;
                when pause_setI4987 =>
                  \$ram_write_request\ <= '0';
                  \$v3536\ := eclat_unit;
                  \$1284_sp\ := eclat_add(\$v3530\(32 to 47) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(\$1284_sp\));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$711_apply_arg\(92 to 123);
                  state_var5312 <= pause_setI4986;
                when pause_getI5000 =>
                  state_var5312 <= pause_getII5001;
                when pause_getII5001 =>
                  \$5171_v\ := \$ram_value\;
                  \$v3542\ := \$5171_v\ & eclat_sub(\$713_binop_int_arg\(65 to 80) & X"000" & X"1");
                  \$v4999\ := \$713_binop_int_arg\(0 to 31);
                  case \$v4999\ is
                  when X"0000000" & X"0" =>
                    \$1218_res\ := eclat_add(\$713_binop_int_arg\(33 to 63) & \$v3542\(0 to 30));
                    \$713_binop_int_result\ := \$713_binop_int_arg\(139 to 154) & \$1218_res\ & eclat_true & \$v3542\(32 to 47) & \$713_binop_int_arg\(81 to 136) & \$713_binop_int_arg\(137 to 138);
                    \$v8\ := \$713_binop_int_result\;
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when X"0000000" & X"1" =>
                    \$1218_res\ := eclat_sub(\$713_binop_int_arg\(33 to 63) & \$v3542\(0 to 30));
                    \$713_binop_int_result\ := \$713_binop_int_arg\(139 to 154) & \$1218_res\ & eclat_true & \$v3542\(32 to 47) & \$713_binop_int_arg\(81 to 136) & \$713_binop_int_arg\(137 to 138);
                    \$v8\ := \$713_binop_int_result\;
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  when others =>
                    \$1218_res\ := "000"& X"000000" & X"0";
                    \$713_binop_int_result\ := \$713_binop_int_arg\(139 to 154) & \$1218_res\ & eclat_true & \$v3542\(32 to 47) & \$713_binop_int_arg\(81 to 136) & \$713_binop_int_arg\(137 to 138);
                    \$v8\ := \$713_binop_int_result\;
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  end case;
                when pause_getI5003 =>
                  state_var5312 <= pause_getII5004;
                when pause_getII5004 =>
                  \$5173_v\ := \$ram_value\;
                  \$v3545\ := \$5173_v\ & eclat_sub(\$715_binop_compare_arg\(64 to 79) & X"000" & X"1");
                  \$714_compare_id\ := X"00" & X"9";
                  \$714_compare_arg\ := \$715_binop_compare_arg\(0 to 31) & \$715_binop_compare_arg\(32 to 62) & \$v3545\(0 to 30);
                  state_var5312 <= \$714_compare\;
                when pause_getI5006 =>
                  state_var5312 <= pause_getII5007;
                when pause_getI5010 =>
                  state_var5312 <= pause_getII5011;
                when pause_getII5007 =>
                  \$5175_v\ := \$ram_value\;
                  \$v3549\ := \$5175_v\ & eclat_sub(\$1179_sp\ & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3547\(64 to 94),16) & X"000" & X"2") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3549\(0 to 31);
                  state_var5312 <= pause_setI5005;
                when pause_getII5011 =>
                  \$5180_v\ := \$ram_value\;
                  \$v3551\ := \$5180_v\ & eclat_sub(\$716_make_block_n_arg\(16 to 31) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$v3547\(64 to 94),16) & X"000" & X"1") & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3551\(0 to 31);
                  state_var5312 <= pause_setI5009;
                when pause_setI5005 =>
                  \$ram_write_request\ <= '0';
                  \$v3550\ := eclat_unit;
                  \$1180_sp\ := \$v3549\(32 to 47);
                  \$716_make_block_n_result\ := \$716_make_block_n_arg\(0 to 15) & \$v3547\(64 to 95) & \$1180_sp\ & \$v3547\(32 to 63) & \$716_make_block_n_arg\(146 to 153) & \$716_make_block_n_arg\(156 to 171) & \$716_make_block_n_arg\(154 to 155);
                  \$v8\ := \$716_make_block_n_result\;
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_setI5009 =>
                  \$ram_write_request\ <= '0';
                  \$v3552\ := eclat_unit;
                  \$1179_sp\ := \$v3551\(32 to 47);
                  \$v5008\ := ""&\$716_make_block_n_arg\(34);
                  if \$v5008\(0) = '1' then
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$1179_sp\ & X"000" & X"1")));
                    state_var5312 <= pause_getI5006;
                  else
                    \$1180_sp\ := \$1179_sp\;
                    \$716_make_block_n_result\ := \$716_make_block_n_arg\(0 to 15) & \$v3547\(64 to 95) & \$1180_sp\ & \$v3547\(32 to 63) & \$716_make_block_n_arg\(146 to 153) & \$716_make_block_n_arg\(156 to 171) & \$716_make_block_n_arg\(154 to 155);
                    \$v8\ := \$716_make_block_n_result\;
                    \$v1549\ := \$v8\ & eclat_true;
                    result4918 := eclat_unit;
                    rdy4919 := eclat_true;
                    state_var5312 <= compute4920;
                  end if;
                when pause_setI5013 =>
                  \$ram_write_request\ <= '0';
                  \$v3548\ := eclat_unit;
                  \$v5012\ := ""&\$716_make_block_n_arg\(33);
                  if \$v5012\(0) = '1' then
                    \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$716_make_block_n_arg\(16 to 31) & X"000" & X"1")));
                    state_var5312 <= pause_getI5010;
                  else
                    \$1179_sp\ := \$716_make_block_n_arg\(16 to 31);
                    \$v5008\ := ""&\$716_make_block_n_arg\(34);
                    if \$v5008\(0) = '1' then
                      \$ram_ptr\ <= to_integer(unsigned(eclat_sub(\$1179_sp\ & X"000" & X"1")));
                      state_var5312 <= pause_getI5006;
                    else
                      \$1180_sp\ := \$1179_sp\;
                      \$716_make_block_n_result\ := \$716_make_block_n_arg\(0 to 15) & \$v3547\(64 to 95) & \$1180_sp\ & \$v3547\(32 to 63) & \$716_make_block_n_arg\(146 to 153) & \$716_make_block_n_arg\(156 to 171) & \$716_make_block_n_arg\(154 to 155);
                      \$v8\ := \$716_make_block_n_result\;
                      \$v1549\ := \$v8\ & eclat_true;
                      result4918 := eclat_unit;
                      rdy4919 := eclat_true;
                      state_var5312 <= compute4920;
                    end if;
                  end if;
                when pause_getI5015 =>
                  state_var5312 <= pause_getII5016;
                when pause_getII5016 =>
                  \$1152_arg\ := \$code_value\;
                  \$717_branch_if_result\ := eclat_add(\$717_branch_if_arg\(107 to 122) & eclat_resize(\$1152_arg\,16)) & \$717_branch_if_arg\(1 to 32) & \$717_branch_if_arg\(33 to 48) & \$717_branch_if_arg\(49 to 104) & \$717_branch_if_arg\(105 to 106);
                  \$v8\ := \$717_branch_if_result\;
                  \$v1549\ := \$v8\ & eclat_true;
                  result4918 := eclat_unit;
                  rdy4919 := eclat_true;
                  state_var5312 <= compute4920;
                when pause_getI5019 =>
                  state_var5312 <= pause_getII5020;
                when pause_getII5020 =>
                  \$1138\ := \$ram_value\;
                  \$ram_ptr_write\ <= to_integer(unsigned(\$718_loop_push_arg\(0 to 15)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$1138\;
                  state_var5312 <= pause_setI5018;
                when pause_setI5018 =>
                  \$ram_write_request\ <= '0';
                  \$v3555\ := eclat_unit;
                  \$1139_sp\ := eclat_add(\$718_loop_push_arg\(0 to 15) & X"000" & X"1");
                  \$718_loop_push_arg\ := \$1139_sp\ & eclat_add(\$718_loop_push_arg\(16 to 23) & X"0" & X"1") & \$718_loop_push_arg\(24 to 55) & \$718_loop_push_arg\(56 to 63);
                  state_var5312 <= \$718_loop_push\;
                when pause_getI5023 =>
                  state_var5312 <= pause_getII5024;
                when pause_getII5024 =>
                  \$5192_v\ := \$ram_value\;
                  \$v3558\ := \$5192_v\ & eclat_sub(\$720_w_arg\(8 to 23) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$720_w_arg\(24 to 54),16) & eclat_resize(eclat_add(\$720_w_arg\(0 to 7) & X"0" & X"2"),16)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3558\(0 to 31);
                  state_var5312 <= pause_setI5022;
                when pause_setI5022 =>
                  \$ram_write_request\ <= '0';
                  \$v3559\ := eclat_unit;
                  \$720_w_arg\ := eclat_add(\$720_w_arg\(0 to 7) & X"0" & X"1") & \$v3558\(32 to 47) & \$720_w_arg\(24 to 55) & \$720_w_arg\(56 to 63);
                  state_var5312 <= \$720_w\;
                when pause_getI5027 =>
                  state_var5312 <= pause_getII5028;
                when pause_getII5028 =>
                  \$1104\ := \$ram_value\;
                  \$1101\ := eclat_sub(\$721_w_arg\(48 to 63) & \$721_w_arg\(0 to 15)) & \$1104\;
                  \$ram_ptr_write\ <= to_integer(unsigned(\$1101\(0 to 15)));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$1101\(16 to 47);
                  state_var5312 <= pause_setI5026;
                when pause_setI5026 =>
                  \$ram_write_request\ <= '0';
                  \$v3561\ := eclat_unit;
                  \$721_w_arg\ := eclat_add(\$721_w_arg\(0 to 15) & X"000" & X"1") & \$721_w_arg\(16 to 31) & \$721_w_arg\(32 to 47) & \$721_w_arg\(48 to 63);
                  state_var5312 <= \$721_w\;
                when pause_getI5031 =>
                  state_var5312 <= pause_getII5032;
                when pause_getII5032 =>
                  \$5197_v\ := \$ram_value\;
                  \$v3563\ := \$5197_v\ & eclat_sub(\$722_fill_arg\(16 to 31) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$722_fill_arg\(48 to 78),16) & \$722_fill_arg\(0 to 15)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3563\(0 to 31);
                  state_var5312 <= pause_setI5030;
                when pause_setI5030 =>
                  \$ram_write_request\ <= '0';
                  \$v3564\ := eclat_unit;
                  \$722_fill_arg\ := eclat_add(\$722_fill_arg\(0 to 15) & X"000" & X"1") & \$v3563\(32 to 47) & \$722_fill_arg\(32 to 47) & \$722_fill_arg\(48 to 79);
                  state_var5312 <= \$722_fill\;
                when pause_getI5035 =>
                  state_var5312 <= pause_getII5036;
                when pause_getII5036 =>
                  \$5202_v\ := \$ram_value\;
                  \$v3566\ := \$5202_v\ & eclat_sub(\$723_fill_arg\(16 to 31) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$723_fill_arg\(48 to 78),16) & \$723_fill_arg\(0 to 15)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3566\(0 to 31);
                  state_var5312 <= pause_setI5034;
                when pause_setI5034 =>
                  \$ram_write_request\ <= '0';
                  \$v3567\ := eclat_unit;
                  \$723_fill_arg\ := eclat_add(\$723_fill_arg\(0 to 15) & X"000" & X"1") & \$v3566\(32 to 47) & \$723_fill_arg\(32 to 47) & \$723_fill_arg\(48 to 79);
                  state_var5312 <= \$723_fill\;
                when pause_getI5039 =>
                  state_var5312 <= pause_getII5040;
                when pause_getII5040 =>
                  \$5207_v\ := \$ram_value\;
                  \$v3569\ := \$5207_v\ & eclat_sub(\$724_w0_arg\(16 to 31) & X"000" & X"1");
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$724_w0_arg\(48 to 78),16) & eclat_sub(eclat_add(\$724_w0_arg\(0 to 15) & eclat_mult(X"000" & X"2" & \$724_w0_arg\(80 to 95))) & X"000" & X"1")) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$v3569\(0 to 31);
                  state_var5312 <= pause_setI5038;
                when pause_setI5038 =>
                  \$ram_write_request\ <= '0';
                  \$v3570\ := eclat_unit;
                  \$724_w0_arg\ := eclat_add(\$724_w0_arg\(0 to 15) & X"000" & X"1") & \$v3569\(32 to 47) & \$724_w0_arg\(32 to 47) & \$724_w0_arg\(48 to 79) & \$724_w0_arg\(80 to 95);
                  state_var5312 <= \$724_w0\;
                when pause_getI5043 =>
                  state_var5312 <= pause_getII5044;
                when pause_getII5044 =>
                  \$1055\ := \$code_value\;
                  \$1052\ := \$725_w1_arg\(16 to 47) & eclat_mult(X"000" & X"2" & \$725_w1_arg\(0 to 15)) & eclat_resize(eclat_add(\$725_w1_arg\(64 to 79) & eclat_resize(\$1055\,16)),31) & eclat_true;
                  \$ram_ptr_write\ <= to_integer(unsigned(eclat_add(eclat_add(eclat_resize(\$1052\(0 to 30),16) & \$1052\(32 to 47)) & X"000" & X"1")));
                  \$ram_write_request\ <= '1';
                  \$ram_write\ <= \$1052\(48 to 79);
                  state_var5312 <= pause_setI5042;
                when pause_setI5042 =>
                  \$ram_write_request\ <= '0';
                  \$v3573\ := eclat_unit;
                  \$725_w1_arg\ := eclat_add(\$725_w1_arg\(0 to 15) & X"000" & X"1") & \$725_w1_arg\(16 to 47) & \$725_w1_arg\(48 to 63) & \$725_w1_arg\(64 to 79) & \$725_w1_arg\(80 to 95) & \$725_w1_arg\(96 to 103);
                  state_var5312 <= \$725_w1\;
                when pause_setI5045 =>
                  \$ram_write_request\ <= '0';
                  \$v3572\ := eclat_unit;
                  \$code_ptr\ <= to_integer(unsigned(eclat_add(\$725_w1_arg\(80 to 95) & \$725_w1_arg\(0 to 15))));
                  state_var5312 <= pause_getI5043;
                when pause_setI5047 =>
                  \$ram_write_request\ <= '0';
                  \$v3575\ := eclat_unit;
                  \$1038_sp\ := eclat_add(\$726_w3_arg\(16 to 31) & X"000" & X"1");
                  \$726_w3_arg\ := eclat_add(\$726_w3_arg\(0 to 15) & X"000" & X"1") & \$1038_sp\ & \$726_w3_arg\(32 to 63) & \$726_w3_arg\(64 to 79);
                  state_var5312 <= \$726_w3\;
                when compute4920 =>
                  rdy4919 := eclat_false;
                  \$v1549\ := \$v1545\(0 to 121) & eclat_false;
                  \$v3576\ := eclat_unit;
                  eclat_print_string(of_string("pc:"));
                  
                  eclat_print_int(\$v1545\(0 to 15));
                  
                  eclat_print_string(of_string("|acc:"));
                  
                  eclat_print_int(\$v1545\(16 to 46));
                  
                  eclat_print_string(of_string("<"));
                  
                  \$v5304\ := ""&\$v1545\(47);
                  if \$v5304\(0) = '1' then
                    eclat_print_string(of_string("int"));
                    
                    eclat_print_string(of_string(">"));
                    
                    eclat_print_string(of_string("|sp:"));
                    
                    eclat_print_int(\$v1545\(48 to 63));
                    
                    eclat_print_string(of_string("|env:"));
                    
                    eclat_print_int(\$v1545\(64 to 94));
                    
                    eclat_print_string(of_string("<"));
                    
                    \$v5303\ := ""&\$v1545\(95);
                    if \$v5303\(0) = '1' then
                      eclat_print_string(of_string("int"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$code_ptr\ <= to_integer(unsigned(\$v1545\(0 to 15)));
                      state_var5312 <= pause_getI5301;
                    else
                      eclat_print_string(of_string("ptr"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$code_ptr\ <= to_integer(unsigned(\$v1545\(0 to 15)));
                      state_var5312 <= pause_getI5301;
                    end if;
                  else
                    eclat_print_string(of_string("ptr"));
                    
                    eclat_print_string(of_string(">"));
                    
                    eclat_print_string(of_string("|sp:"));
                    
                    eclat_print_int(\$v1545\(48 to 63));
                    
                    eclat_print_string(of_string("|env:"));
                    
                    eclat_print_int(\$v1545\(64 to 94));
                    
                    eclat_print_string(of_string("<"));
                    
                    \$v5303\ := ""&\$v1545\(95);
                    if \$v5303\(0) = '1' then
                      eclat_print_string(of_string("int"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$code_ptr\ <= to_integer(unsigned(\$v1545\(0 to 15)));
                      state_var5312 <= pause_getI5301;
                    else
                      eclat_print_string(of_string("ptr"));
                      
                      eclat_print_string(of_string(">"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$code_ptr\ <= to_integer(unsigned(\$v1545\(0 to 15)));
                      state_var5312 <= pause_getI5301;
                    end if;
                  end if;
                end case;
                \$v1821\ := result4918;
                \$v1820\ := \$v1549\;
                \$v232\ := \$v1820\(0 to 121) & ""&\$v1820\(122);
                \$v1545\ := \$v232\;
                \$v1818\ := eclat_unit;
                \$v1814\ := \$v1545\;
                \$v3417\ := ""&\$v1814\(120);
                if \$v3417\(0) = '1' then
                  \$v3416\ := eclat_true;
                  if \$v3416\(0) = '1' then
                    eclat_print_string(of_string("cycle:"));
                    
                    eclat_print_int(\$556_cy\);
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$547_o\ := eclat_false & eclat_true & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false;
                    \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                    \$v1527\ := \$v495\;
                    \$v1810\ := eclat_unit;
                    \$v1809\ := \$v1527\;
                    \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                    result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                    rdy1858 := eclat_true;
                    case compute1859_id is
                    when others =>
                      
                    end case;
                  else
                    \$v1815\ := eclat_unit;
                    \$547_o\ := eclat_false & eclat_true & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false;
                    \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                    \$v1527\ := \$v495\;
                    \$v1810\ := eclat_unit;
                    \$v1809\ := \$v1527\;
                    \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                    result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                    rdy1858 := eclat_true;
                    case compute1859_id is
                    when others =>
                      
                    end case;
                  end if;
                else
                  \$547_o\ := eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_false;
                  \$v495\ := ""&\$v1814\(120) & ""&\$v1814\(122) & ""&\$v1527\(2) & \$547_o\;
                  \$v1527\ := \$v495\;
                  \$v1810\ := eclat_unit;
                  \$v1809\ := \$v1527\;
                  \$v1808\ := ""&\$v1809\(0) & eclat_not(""&\$v1809\(1)) & \$v1809\(3 to 10);
                  result1857 := eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & eclat_false & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9) & \$v1808\(2 to 9);
                  rdy1858 := eclat_true;
                  case compute1859_id is
                  when others =>
                    
                  end case;
                end if;
              end if;
            end if;
          end case;
          
          result <= result1857;
          rdy <= rdy1858;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
